`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hH+7Of7V0HrZN7akhr/PGWzFYMFZ/Rw1Y0MdJHcXbDfy25bCrbSAgiAHzjAOItzVH0GJHC0TwaAh
l8lQ6Djj5A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AmHoZR7VmEL3tVmWsOV6IVQew/VOu2KAm4f6KJfAzXGRTTxsXlPXI5eOmXy0OQc+dTQXlc4Nyebk
WOd+g7avEM/H0dDmrnyrAy4xkmGgWvy/yoSRg2NcrorlzU30DXGyLUL7cC0fGGT3+aYDfpalxOxG
vMlnYmB3ol3sAa02k/0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quTe40cgTFzwGZ4hh0czXTRPjRM65yQ2xuoMk4KWhGRBXqG0mDC0qybq0KDkzMvHMO9o13XXh86J
3lmXd5z2U8qbCCQTiQ5D5fs/vDyxOt2D8yzeP9Nz3v9pLob1z25U2A3IDkfdMys+0lSQ2Kic2K7X
M9l4gP8XjJ7XaZMV90LT+K3emy6GtwfHL1RmLLmz0wvq+4goCsSl98hEr1onaBQ9FjjXJSgHTEoZ
asLa6XQpuzHvUdrr7uow2fs6n/v6lPMa2QIEVAOBRHRZfcfQ8mCrRActebecw4kgaKOLxGzIWyFi
VJjLlE6Keg/yDxLLEGAzIe0fXmz5IeT0hi9g5Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e0IXUCRiGRcDhitPNE5pcnOQjcFm6XyOGSyf5ehAs8DfcUjdAyC39hcyh7lelM2n1wk5DOyQUYdV
sH1HD1x890dqy0Bm+/WUTKfxQ5I0MfCdzTLMWpdnX0TYkOpM7Yw8f7rYC6qJM3409nB55jo5jbXs
BAEUxqIp85fdzNw1bsDtj4/QyVBwF3hP7nFhpQv+EKdvqv8Q0w3KT9MgfmK+tlzpA7nQq1DUqyYL
tY84oCcSfcuA/mVkkAZzSZD+v/Q3sdnagb4fc0bpcJT5TQnRzdluhqgGQtVo9Hv3B/rAkJ133atf
AhgpSKBM/HuMkZ/NgBMJ7PD7eVL6yIU2qjgBTw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h5kgqPrm/ghas5o50sQF7CkRrd0UW9+3Bgyf9II/ObYHKU5WTqvdQVx37RiV6Zuwx7jY8BKGUrC1
6GljDBL3LJhoaR694OorSigRqGQq9DlbWwvPpubN73/pUcAA/BmXyPJ11iAur9DDz8dL8u0AIVBZ
JMEcSp98XKgEOnXtjaU55MTSv0JNClbz/1GbpUB/la5GmUUPVd9VERL915SygcAxXa4efzVDfNQe
TDR9Cg+V+hNwUsZ4AL0NwCpeNAD+IBeM7wr73ySKSUjSInxlA30lGKpFr4nZ6c/01uzl+nrIAdot
iHHtG6uFhJXK84C4UUrX6PN4AXNBi1ScXRAvVg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qMPgyiJBLpyBHm6njnuRl+5NmZjHACVWOf0ME8HZlaAMEUuZ00geWO2DJ0BCcg6vVw2jNUSHe2YL
wAuBLQt46RfOun3ifJd0vZ0OhmxMdGpmaBkF+pDreoI/Y+6zbpN9NLfWQkPSbXW405FftA6mC0LY
RxeVKPNt7taRM3Dn7tk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GOYJBmvSniPrLCFEvUHh6c8XRUg3Opfv+CEOXcm6o+imohXua80ifxh90luGWez6hJmfSTaDELfP
EFF5QnNkriODMphgc0hRiy06hmsvCugkY/+lnM1+vmLXcLsYksCkRp1yvno838j5TK13b7OUrqjF
fpYN4rWrOt+Od0qedbEyjVw1DaVbqvMeSEy09YrquzpAB1Gn42zQnRqbZyB3P7UxKxd6Je78SneY
ZTMyCwaU8UpZ4qBnHHuRlhiw5mnZoM9BogaBHysLvo7BZaDOif/Zebq6qPrmHuj0Z7B8J4XLLpKP
kYrrZxtmMkKcHsR8kM8j5XlIL2/TVXXoecYL8g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QmPcEzlUpwA8HkI5E7k3BJ8/+g51Sr0bTjftiABHZ12feKb0yyUwc3DGo4XhaK2hwP9A/eEaRoma
DGsRKeLWw0e3ct2vRi8ep6WFdF7j/Iem/cY4NZlDwWOsU5p/5aUY6JIjthh9yRXtopvvMjCYzfsJ
/aV9biiKpCoceP7BX9BA/fsNJMkN6Uz53KSeUPzAHhAjmqbPrq1tftbyHQAdeTBIITSgKrbeoJwD
MluQlsoQv6FFc/AG8Xo3Jw0Xz2SIjACi5gXO0Om2I4nU923OlhwwBiwNqVm2ItyIp8VbqOkoT31n
b3utr1501a+m4vRbYf1P+coW4adHWojl7PGtnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 59568)
`protect data_block
iDYfqNwlpRopY+1YWynzvdDiz4ihvWKObGnB/CbpM0ndy3b8HYKHOYVxW73eYKS8P37UZXFbZaRn
OswUg1hlZrPhTv+I3noV7716GA6XzOsL1/Hbb8a/r+QSTiBjM1cmvaYBNGTX/ilxwz31H4+MFg++
vcq2XisUuKeE7zUaJWwseBe5MQAWLLNEtUhWoMZpF49b4CcQnEdAnTKcLB496iJuvLUwVVAi0ukd
nhN8ZnoLUX9oEXL73zGifM6DmY3OyfhQ60hHh1oZm3W/Sd4nO8l9Hr3YFDBAA1BRQ2Nl/5fJrY5F
kU9ywHSzs63WxSAeLxt0q6FLaCBKPaD8mjGsnojLimL4FqUIpUkqTf4dfhEyU4EhsDq3o5o483gb
zWQe5N0GYEbQ/R1nDF+y+8XM6al2/FU1bTYabfuOPO9CcMFaHgLZ8FwuqefnbtHurbGjWPXLNmo2
jL6bDTDLc4XzPgg45t6pMYCQGrdVfNUum9mRCPrbbbKOnk4PjfsWGIWnSCGY7EKIiapWaTTu7iDE
DLRAthE20jgOVj6YKcVW0n7z6h4cR5bxmL3muCNcynWTYQK6Ak7UCIQSA1YhYSogeMpAO8iu85cL
VRfY83NVzCkYCs00jm091QgZ5XmBejFLDsPE4WL9wpdZubOhAdTWiJvGqlxVfkYXgQQo7ENItkmi
RtPWxu4D1Le6Qp0ttE1LjiP+RDcHZYY5/geSwziiBo1EdsUEjX2pI+8TrYle4OBJiSJI3GHe2eeE
Q+8LK2yW0AlIJa/8xwDun8/eoyJ84roPG/UbpaNMOFnZzjpS4Lkr/LOtqv7sSRPaLX20iXms8bH+
RGR4S5rPDTDg3N+gXc6rjFbEAMbwu0YtGk32m/8PyZHf4XusjuPLmNqOThVcvOvYp16wHyRsNIiw
q6aG2kcyVlriJ8dwFdkyEjx/7biUfrPFLP42puSJ3vD3b1zj/u3RGYHDyn+QrMqZBZAwTQti+84x
sVlaysFGZ6tXVOemm8LWLhLaTrM4/t0pZ531qgbkQDkd0RNVFsKm7kUGKcP5WB1diudBD4TTnond
F+tf5cNbdGz8PWjJdFtjtAbmqA13Ouv+SKw4cuHOEUgYP83vYbFVX29eDOF0v/ZzYYc0yPbd+8cX
3TJR6AOxIIbWckj0E+2nBOTNRLHq8ID8q6L9eWETEGsWb0AKRVjddK5OtDDVi3McDhKWvmCyzZy4
Prdwh1XXISqb68GsaU4tXPPWDLa1T0UCggA7rQNWpwld5xC2E7qwR+z/i6xfosW3HAKZ+tLwfhBf
aU8OlxBJg0ci6IefP0fqf517Z5bRe/uqk1fNVI6k1WWn8TOGUMhDZLMxcfUTYK83SOl7IWi/XcHL
FwWLv3sIu130nCRPko3oDw4/O+JKGK8Z7wYgtbraI43VCJOug9p9tNbhlqikEE03jKcrdqt+phb/
PGjZiPcHol3gTF8UJMGntN/L7WU+8+2NqPAII+LES8hqv1b6ITQ1cXsUcOJMvYNtKOagWeySQXHu
N2jQ9tK6KLZVbaJEKB/vxVyXdlLvr/Up/qJKDWMQoYw01VL41Q/zQ6U9LFEwg3o/eDEyzW2SfybS
SySzONUxVStAxcQMNHRG+L1gwFadBPI6MBQ8xkyd3dN3mSA7L3d4KSpyQv3as9xa0e0l8/fo+jHL
HJRnyvDe5i6SLIg/y4Rt06XdzwnrhGAIDHaEQmVFBvSK1b6blKSlPe+PoZXoizHidXYYIm4fDNUe
qLdGDoisCPjXy09PDSkJ3VV0ZjaL/ZWJYoi861sPZSI2RPM1cbRq4YNdiwVbD+fsSuwXXIj+xkp6
w6VKPuGiGtQK0GLuPg2nDZYXh64H5MmLI43qlU1kSaE38S3XyOBiJiA6h1fCxLjSFDdgUmsAhi4/
CBxf9V5LgVri/MZUzQFS9JjxWPk1vNBAQ/+b4SbJehio3G2ouewkWLx1pUQNKR6vfZ8ZOjUKxPpw
NG8GEpwbr/AEUWzZpu+2SZhobiE2uhk8CEOwmV5i5F3tmi957nOXK0EkXDau4cFSlGODrCWQOpuI
depvSK22KltcbZ8Wvqhok5dHeDe3yjB/leGQJo59L9kJm6pq/+h20UzD8L5D13ZexwV9uK/IC0iy
DSpVze1IWzg70tyNVORIJ01//EeCfXXf+IoaPdPmkDZJrVdH/ce3EN3bvRDCORtNIzzD2TwW90/v
+SDjNJSNpdG55vLBo7xLYyOppEBgxKCQwOulA0t88pSrQQz4O5+uI7xF5/EIoJITBGWeJvN9ru3U
Bvq0ZS/3rVdDg5QwG2KMYHz3TpRCrfxSsEADu0Ke5PUoG7l8sp2CZkXrz0nCMfEBpbYD3wOPXNLc
ZwDp+jw5SXtL48Vi1GqPO9swRDG3v1WEo7j3hzmUWbDmx0Uy5nXj99EYZVWkYDSCLoVV2l3p+ieq
o8EvsFB3ifI/bbigPiOawwy6pG4oTSAlIk+htXgCZwg3mlqR/7ZV9AQAk9uBoC86ODi1dNqkvpdI
EbfgNrBxiuoDpNrI2ojLsWbeHFHt1GQQGh9DsWn6Sn8MtrzpBEJaFrkSRUPjylMePoKzNPE6GIU7
HY/yq5TUbhV1WrGroh8rDsy3hEoXy2+6FyLRRPCACi3YqMs8zLljTmR26Q1sELa2deZRq3TlyWEG
1VXXLXLWtCY2RmqwPTM8E/3MILo6PoiitjV5iesaipnwIGTe1XrU3ZYhxY9Rnymm9tj5EGpO1ke/
yc2ExZEsBrHGfN8t/0NCIPQDpeA8jF3KRtfOpEP5wwW/tr/vF+HbQsz5BGcD5tOf/FFkXXF6B6Ei
BoUenWX5/Vahl0MgrgVix2BR2ZIdNU6Q3HtjmirtcPMrEdmHmWdnb+U1CxZyNg9lNIh4cC6aNfSC
t20OSirGEuR3u2/rW4IIe4s/JsGqiyMTR33NyCI7fEpZIie27TwtX1QfN3Qyq7MfQMkkmqiR7gzF
FrmioXk7GflyLO1q1i55kLSUqOsfoqWxu9PrOUgApRCZzdOEGK/fRGIhLZ4QEvt5vXMyE3feJwgy
fQevwHTLDFV1THHE+mrHnP0p367nXNTRVY4km962bYAc7qjxmWWHgBbZ2hOU87P5LHUxMkfvnCyR
a2NnZZXHsMOfavb27E5bR3CTYIw0l8Q1c7P9XM1NPdnKdeAy6qGoui7N+8ioFE2VuwMfAF1Rafic
RdqEIXP3Zrho+8dm6mXhQvLhha3vH8MbYhhemKHQFhwDDE7477iTWlXNup+yPdX8hL8wUq2dspx3
zxWTFR5hp667ZuIHx/LT4JjscyzqxLl6o2tJniks8AUpRbUWJ/JMtvrFzbitF/C72YSrSlFMlEEj
t2Way/8FRy32hqYxRBRpsm9NmlmaZFDcmB2dBWovVh+MnWaqnqA+CI8BdJNF4fNqaaudSLSTlzXA
0KSe2YKYVAtqyN7ulwqtX5u0rWbz2BCPXuwIOBmcbWzmtGRZTy1W47eYEw/NBQxFgFPkZ1kbe+bz
lCP4eIfn+rUZ8L7GjVBmS46GBIE/i++kvuJDmyqXRm51vbSdQK6tWIBfb5luuHQ/2DuBKMgXZp/2
R5rID4ot4ImnHea1/UBfE3bGiO8Bu4c7DH9Tuyh8mFFxe/cr4CIzmjHXWjMlcYOR30p4vW+AP4F5
UzJMRzXkaHfmWk0Nbdtv9pZYW2LgWcQ11fNGPiVNxEI2x5057PQqbz3yjQOpmLYOB9A7MBJBOwGj
s2XXdN5aMQaLFy4mu9FHuVhBfzC2rPT05UGYdsixQlAKHy0ZRzQ43cf0zKXO6Wlsg+cWrG/o7jbM
b2YMXDWU+Abp3WUc7BCX/TLoWaxKFU012xpcReDz6UFOEnInofyh7D4d9lsHa6SfJ5kH+7YvM00B
rRj91v2dYIvAEtEHhFRxmEoOrkmVEOEtI3ZbvKUTky/4eGFe8FPnrnSRYySNYbxdZZVcstHK5b5h
BmWScHLNvUjK8WeHTIjThswsey5PSrIOeuvEJDF1LKQCSnYV9fsZj/pBhcak3eGtYHkG6U2QW9OX
EOlr2wuM6RN/Ta9h4WWTDSMiR9UHSqo4p+SEWxwieCggM8EgtOXZrA+r07JSWFG/NFO05hJT84xR
7VQ7luYkV9QBvs7X3kx9k+DhFAvfr0gGHweUY05Z/Xxd9JIZsLr8Dmmk3vBv87or4SM3KabSEkgY
klLZnanT8XRb+Ojnvlwa/PN+ipaiqHy68BJ7bq97TV8+NfRGET8p7qRPAsEPeeGvCy5Hi7p7SPXM
Bb6zK2pftwPDF5Dg9ZUaAI55X8yXq4yY6lsIGiWWtSCU8LEO5+6LZBan7ml5O7z8CsW6L9/j4N/M
Nr+RaBUkMEC3Bfx7IGQOlBsSgKCaYwdOan4M2mzezJs0iR6mVFxR1epcAMywR4zBUiVt8bLLTqhx
n+NRabJ5vkqeYwbvxP2yYDqLbu+nwbeqiGBtDQsLuUjCytJNtQe5NqGRP1y2TFaWW75ttRNUCBsz
wVIo193bt/P7pDPKneUWeQnfhDPfK6kbZISel0L4YkLm52l/e8XyR5jWk/mJgYtjCjgK9lkr7Kl9
pcDB9pbGI5Eg4sbxfCTwkdO1iB5+uw/MEP4dlJpIwWSo+467JcgpDd8yfrm03AcA0kJLJGDE9yvs
eDiO+jOYx+AX6CnPbznTdYi0ZHQVIEWCDVrk7LXy0jJc3Xe7XuYkUjUUFqSXPqLwvaf8ZGvCP4N1
71auDwrDQ8Ndd2dLPeAWjT3RiJlhmTNq/prg3esDmWLUmBrPoUudD7PvHC1NsqiOPh2XxSzXiQls
Mv0sth8vBbQJDJpHwb9WE7mUgQuDDz8UFeLN7+5gaPxGqemIlLTs4zrBvWUU0a8iMIf5q5UKxL53
1G2/iU0YUs59mej63fNpS2ee/vaN8SCgzS0AE3ASRTHdMZdHkJaSZ8/gYPz5ZFOY9GGZVjoFGuoM
aoVQRJaQZBpmq+CwzoPAjeCCjV2rkrJRONyd0o1TGL5a4YbTvwODLW5cuRzbTID0mm0EB3XVumrs
ofFqmRkauwS7lu+pdjyrRTDn6cdXktgI0+UnQTy3wMm1y+IVkPQEhiy8fQ3KBUQ1vp4ShjafffCa
N00v2Ce2JCYLTpZJTiEG7uDuPH/XN3/OU0MghGj0NKl5zU+SAIu3PBiklYQ/C5nZtJfVoJ2UjTiv
R/UaykvKQXKmBG4pXsggcJGHmpxpm/sVM7blumkCmvVZ12devRgYmMD022tKmyKNcFmMvnaVLNvK
PsvhYep7qEQVM7ZnldLk7/+ta0rzLH0lR9ZTeZYwNtK3q1Ei1AlGmezKkVUMRj51ELYrFgMtv2Vq
A0ofocwP0kHvM6334r1nSDYI11tKhAI7z1zjL5JQRF2Z8MnGd4mkpVjw1HnQBNteHUcbIKUoXo1e
gYGmcL8qwAbrk5UcwyaFwDGDhtQ8ErQBhjyv31H0IGWb4l07MZ3drYINlM8zqDjp/r0hjQRhjwVp
4q3N0X4/0R6+vqVDJhs69AxVlXcotGhB1/ukgqBh38XRmwx6KaoVbWrfyhnb7wKSRfEkGRyyClK7
Bm7S7Cpq4BtkwBqnSYc4bY+/EwT8M/+3To7y0/TN3dTGINr9F44Li0utoEM8U8LNJtMT8CoAiwQx
bBYrfa6IWwm7wx+2Fnq3AVlZ8bjXyJ8D6zUDRJYoBbU4ZyTT8svlYuRuf0TYUVF4hRzdFXypB8AR
JWZU08a+OT9sXx+Xw8eXvZ9zuEYpyqu6g+WwnyZJSEqLlGXn0QFH0Z2gHO8zjIdGLWZlVUd4pAFt
Rc+bbWm+IkgZEbuuuw2yji1DlWsAc6PlFfefQNpzf2a0C0B0SfTyJU1mhkePZixZ9YyGNWkQJyVn
jQrl44u35WUyO6iY7iSNYJyEJBo+CEZqiaW8f4S1qaqyshZz3TbvPlG5LXJc7wn/ITgxuGfa3Xe+
HZlA9vGmKb+8jOWd1O8v6jsUykI0/jw/efOdR0Xydk8swBsY3asWe2GuwneF0q9vguKBCjHxMyT2
aSvgGuUP6bNN0FzkxdaO+kIv1Zb//cqunkA+rRUwbx5H5HhhwddhoZw+RtsiYBEC7l79cWeebMuH
1FnVOYUtbGc+X88Agbp5+AE463lkJOtzptBVOX5dQPDgYmK0SgkPBxUPveTOSN6XThLaH+OG1EIN
CwKKbf+0fh2RTVdVNpl1K1ivVqXb3srqXFQVXrl5Ct2OwdVXXeAHEkKLaTxOGQ43tNfdORLFgKoU
uiZv9GTPivxK+U1XDhegkLYSvcc1Q1u1qrECPts11JK6pUwoDpNGzgQCgBIU0OiqwqbLbC40Im71
Vk53exUaeCiFBeVQP1RrpUby3asb4yToECcYo0nYgedlEnbrR8iWCj+F7lAyEiQK/n7yPHvUQYJF
Npu0m+3UoDXA2RctzRKhptPs06fqv8YJh5MwjWo/1UL8J28V2z1lhTiGxSz6afoCk5FOqfnuYdl1
n76Bo1yPNwZYUsxvztIxRwglnkuQ7DvJsT7D1vWkvbmVOza7LDBuu2z/U6v34AeyogoxvFgBMz+u
445FXhfxo/WiddqXIj9uT3U/WBX8pSxdmpI2EpGj+31kuCp5PwXb4kDAwky3k9zabGknKNvuUYl8
Lh3fH1zq7jpQiR+dkM117cLXpAECQSkszstPzA1dv4SylsNNM4OHmpR/50cRQR48Fxf4p60vzRvQ
bRoXxReLrHPf9akR0MnEC9XSH0or9oBDpRHOEgNfZbvbhyHYIArAT5KPA6Fapzwt9nSIHI21h53Y
hLAlCoqCaUsuQJxd5DyCYtMk5vx7SniEnhbMzBy4xT5TLf8ZWWyKG9oeXRd8DFnMlzwA2IHyONMF
nLk446Ns3vnFtSAC+5n2ZUdZ4+JST07r4GmhfPmE3VNXyxfbuqQ9Whxl2E/N8FfMIgsrqPCPNL4J
NNvvtq0a2mtvMvdNuWgn49RIJK2JkI9kD6b97xmoU1u/GoMueuZx6DEHyYuTOXgw+GssrJEm9bDp
OstFyknHB9hgqBeKiClXhJEWu2/lCihVBJuqi7Ezrc+JiCxrJJBQXFH+8JO6sWP51chcFfXc9szM
J+fLQmbxBnY7/nou0TcPazZDFwyMipw/4iPE1/SMX11TELRsprLc+ZCV0Z01DPPYvHRcIPoSlzrc
MHv4szzY+XynNROXDUYnS+zp12X0Ci8lrlp6dLISjKyCK6wEEblVaWDMTb0Wf9wXh6KSglA2470u
jj9U4qK3vIRrY3E/jMc5w4cnQxLClSZZ5RgD62Gj7kzwrrizYGOoYuM5s+X7JxUvtEmBN0Mz2dqj
cTO7WVaiy9k13ovEc0G9Iao+lyNuhniBYiogBRdqpp56t7V7pD/NEK11fSbNcasgCT1QOPjcP6yy
5XUT/orJNghN8tLV9/1qHlB6vWbG48RPRI4Sua8ui6ilpXili0CzNjaNu05/uZ6NC2JRoIQ0rvlI
ESqDa0J5n8zGwq7/1gz2WxJahcLP360I/Ua+EopSpE+IhlJqcBj2dSltO/yFPyYGZBn/z47mbFP5
QMO1zjAWXqjKzLjjJq08AUzaQRiCWnfi3FZUzA8cRGjTXPxAqRZW03HQO4141gzKo9GiqzM3QaBu
XoBDiF5gx5soX/wy9U/Mb1eCt8DKR0m7qoBwUyJ9FbVGqcRKMMsmA2QNfDgYbfrMw5hGrGLjf/c4
/k+x7na6p9BcSrAE5+y3/iXWo5etRIjH9zSXME83xSGEV6bUxyxn9HuCl8qvuFflY4jtbiUCLv/U
ymnZGKUCe0b3i90YIALIC8JAdY80hrlbAbkGEqgA5pqmchB6IdcA7xo4vY+bkvzkY6O/4EaENjGH
gHCWJ7Zv44HJqyz1UljbHS5c5qV2iZXKj+jjpmMB6E/fUd2YZXqp6ZEPqETKIGDTm3MOutdKjRxY
pVTiVcnPdSAFiohX3LFWyNVXheK0dvTql7dTxiHkbVZc610YSK7kcYTSeKWNK8UczHNtx9ai4ZtF
DKjmbGtAXhlIUFxdVhrsjGruwNsT1el3Wn0S/ma1C3sK9/Cg+Vuf3IrMyqaCXNAZYZyBXYgg2fzs
B6k2xnyd9A86LmLwqIcD1MZ9AKjTnTa19SsKEf4FDr6Q3dDxcZfQTmF2OYQJedR/KCXQ4MFd0VxR
2EgV4ts+1A4aSxz+ws0SRU0G75CipM4Ylxgtk0gfzLhzNqr6+zQGD4kZLohMDNRnZ4gA1K9tBf+4
qgEj0w0Jg0Ga+kXuFvm2FWoYdkJdpKsp3Nzuw6K31WzjvlgF6759rSZZT7VzpoCpUQOfOnWPjzYT
GbdvN3xl3MVKWUvzQYkLIczzHdh7jwHYZslwpKA+HFicKCBchu46rRJCGOfSlT+3hEgx3ZlwedXk
Sab4kpsiIyYH//jbM+0E7AfnnNcUXkFwVBxhmnN6ZNQ3RkAYrRr7YK5ai+ajsfK/F95LOq1aVaXb
tCGZMBoIiGeb3OyUldGsvmP2pgpA+6/VyzfCeG6lRFGhbczqEvhgTUAOs5q89W+fP+N1kvMB2RVV
vfFpIrupfNNzJMlzb1Geb/k4QROKVsDAZ30fC5DhLVDpqB1KQhePh240/qLQN7CZYLM6xClfOXpH
Cu/FeeE7Uc3z/0Q+OqnF2tLPycb8ahQsmRVuk3BG79ox705wbQuE9iae9y85U4c27SNjRYpamJI7
75jt03XjNQTZorUPaMeHzxhx6EMGOO22/GKeN+pkUY9WXFuVhndKE5Wm5HjbNJ9NH+aDU9HbxGFs
1yfWmKqKPdvG7WtwrYA3outvxqmPszeIjTMdcOlzAI190n3OnNhYAcCJCDfAPNud6aJms5Y3rw4p
2Wx+sOf8Xu2BmofffLiVvTvbGYvvOL0boLxkLc2lr56Fh57m3EcExHfvB8sIXxpoJUcCQeRhAXQB
PQTd3MpZ48snw+DMRJohp3iVgx0QG0+Jy+k3kc9IjG7SYhZ0P+M8Q/P8R5j0GLktw48QHcZVrbA/
zq0af0iTsmmGnYDiGfcF4htBjm3zggwjSAJa87ynoLQxVSJCCg07n/K8VG5oEj0WKnSBLx6telAZ
c+PNv9OEpdw/bDpcqV0KnF2+caQcVAQns9q+2q0hCEVwA2ctK7WTCr0l9YtKAqixcONXwwslO7jC
tyYI6XdonrkyMUH8S5wsZSyqL0KR6zx3QlCUPerZffof/0Z8S+rZ35oPlNmv9zQVIUIQzhc3jusI
BQhoauyp5ioYUadHMkhiZMbpHOZIF0Z9JCQaZF8OLk72o321xstcJAYTPgGz6bDHf6JDuzrZcEx2
W5wqW3BjLqlI0ruRvwBRmV1cGFE5UKEdVeT4UfrcH1U4ZNWQe5UNRzAUdpJB8vCQLaF2sC858Iwo
Q0mZwq/ec5YCkW7dwJYZrAmpbUfM2bZ8bw6QGrbjIdON+kgxMyFpzq+dJUXjblQvmZW6+P651c90
LtxpigNsVuTClE1qzyvMGDJ7YW/fDbLMl+uXtFVHEXs9MHMcVEzt4eb+dZ5XMqHeDg+SOz+0PqpP
3SCgBASDyRMk2G/CxutVMoFkOPH0MNy3ApIXBt9rCL8il63oXakS9zNwfbaXCItNVhwafw1iduCD
6MreZyr9/HdByjcN7T46zqLp0PxOJWLjo6N74X9JwjBOZBDCW8SOJ3pZQ7C1UujZor8gxd24sHwT
Ss5uHWoUu/2s4WVbJyaX7fQrNTk/q7oVvo6TBFnwsmHg9leSxrQdJMB8IlOdl3OaxLCbLAJ8vnI+
8D2gyAl+CB54AanpLSDbdrx759U+37V6bkvN6omEm/a4gx6Oy0Dl4uWZvp55VWvO/Cqva+fgaGm4
UDsnaBsUVK6sa0jLMyGOeanDqGHWp5xHnk+zgKM+fzyr9Eywa0FCozH3NKkuFaEUPQSKPZ8k+B8q
0aky07EAaSu2Xr2lq4dymANckDHCzpv1WOB5PW0a0/XnVdd/SW9J6u9WBhTpkebm1lq8ubwn53QQ
1sEawC8xBUszyUBy8zKDm9S2/j5v1VLpgIiFhJFfJ3o2Zdu3trQgo8x+vwtBnFpYtz83l9Z8Pucl
Ozl8OARE7CzMWowcfWCvmA8eJsJGbG3weLQkD/jwWvrvIZFkLyWxM+p+mEqLbss6KpTa06bq5gNn
6O54nNUK21ZRLwYSN3ITq/17/D4TER0jWVIe8z1qLQcdKgZG5Iijw6JP0Z4D1Hb6ilO9uOzAmNWV
w65sReY/MKTzfX4FigM43fAkh1MJGNGMFDrU1HBAEWwHh30hb0UIKYvn8WBRPPMpNvIgpv45UpR9
k+44KcR7bog8HskhaUja7r34R1v3YRP0I0W4/4V2IMaICI4PZKWlz3uMLGqcfglZ/krH95om3O8e
yLqyPJUl6qypTroG7p//yjKisS94i6V8vS2RIMQ1YnHj1JiUrD4A7bgPd0edFrq0dtVtqitTZuKL
3LzFBEvWbeYeyR/qSwbnP+p0FVd1RdR22iH/pqbzsQLOv/gA7ME36T4RKXWEEz++CVsLCEfc8UCW
qAjuIPt7yurZS2YDMi7LIwClAvgZvvhPxlgSrCIjyndCls5qcwhEWpmQetuYWwR4LM1TgCq75LbT
dDXH9dkhWGIHGIZEQSun+1lU6crYxTXFoL7WMJn8GlG7h7pMRoMyozgghrRoO8aHUfHx4BI2N65r
zPY0cLSGXqm+XVw/1lOPAvL9xpCH3CoG2PtvtiXu446LS7LrEddAQ3k/OStxScT9BHTtXD5IEJqS
O686Zk4H5RgBswOZPdPDPNTtU45Tiagc3v+svD36hjU2419T1YF6qVzhzDf1RqfxmesvVyM3x6IA
TyDXZB+7/mJ2328pj8FpzPbZ7kVOnkvJog78vh6WXdv4JxgLSWfXD+I8j9fJeLn6eoClSw1okLJ2
8CIHB99/v1SWgBJc9+IbCJahe7Bv2JC9+yRoA3wV+J74zpv3w6o+sRTc2cecUsTz2apBZ4OP2N+e
4tDvbFFvZPTRDMyz3n2K26hRmqPZyf3ph5soNYokYBi2jMg2YHNj9cpnPjS+bikXWUB5HQhkOkir
W3/HTLJgDWYvbljtkgcCgFj0ej8SSpwsDvQ4G4eqD9GvQ/zhHZdFAZL19C/eukyb306xZlqnlKSp
tQg6eAb6IrHw7JZEPGHlNDvui5UQqTkGDIJtAYaWlpBllB/qWl1A01uEeA9u3jgjNz053D25MBHV
fJ2e3UC0+DtRgOadjMDQIv8HnA2C5+btiW46JwzmpNEDzjkB7pxrBQfJF9f1+rPnmiUNxT+1w4Z8
JXcWJuD4iHaPNfRmFCu5uXlcvNpDIFaVbG9pprhgQKkvxmE1dpcsvDQLX+27G78DC7cipbb7udUN
aFpc7MQ3WZ9RB+v1InLsaScQ8z4gH4+GYBR1c6WstKxqTQ9De/H2/LYb6QTYxQrYYpOaYDH8DO8o
tr92RHojRdQ0t78L46CIgk5J8ceo/dihAk3xPy9nm1NgC++uwqn4x9l/fEab4FZ55rZTt8AaX/5A
DB4nmTFQpFGTb94R6WhB3kRLm18VrTLiutHIuKpw8n1XG7IPR05TJDEdoNRu1ALv1BrSF1b7Hema
epw9U158CbJe2ZWnguGYSdnBaMwczSkRw5ev6VaKCd6lMxJ61Ns22YVOgshyXT8gWEWW0IutKYiU
cU8jzG2Ib54YGUwzRIIBY1+KSMA2NcSo4+fS6r2rGP6SQ4RV+AP8C+VviUrbtb7xuiPBr1FQA0iE
s/4htVb3DJSjZ649t1tL2TfsV5cea/ICvtwE3weuqgnK2jQd/j47cSdArj7mxFTH6W5CfKlD9FyX
fqb0XEOFSvYQDzgquO+sR/Yy0En4OJWnMbiJzs29J2fz1vMogGbof13XhmqwLD9t1RUYYC5Q1f6f
UyfGV/mMv/hLyBeqajFzjDOp5pTzJ4xmMR2puxwZUrI9lZdIQgdBePK8+hY21D+bt6N998Uizcrb
V8XcHZN71a4aUlTkoP6ugU6aFX3HzGFl6y9rYZS6RxytkO3DQB4E7adlkxcpKVrV6QyDGN/T59rz
0Lbk3wYcm4p6NWwXPZ96vWOR0P32mgseyL4GxnE6EA2lWEoGlvZc5WY/EF3ns0HR7M65x6St/wlj
UaIviDXuYeqRb87oWjJPsXiSTmFd/bbD/7Zzg/wpsGWXuZEVPdukjS/kHvruWcUs12y3CX+YhKNW
GJSVXn/cAcU+6filWr5gIACgbu0AdheZIKbPa2edV8K5YNHEb4rliO2Fb7qVmxwy8Do3McGFEn9T
rv2wn1vp+UDdQtKcR4jZWP+jjBPfSvEbAr/X1eJihJ60ftbd0uba6OR/50VFiCUwdo7M71We7ntk
opDWpYNROxm62OO8iu4MerpKIVbPKE107tNWiUPksZHvNZfzd2EInVkWGx734UMxQ6F8b1e7CyFX
7ZeWWkGG8fql3DmJjbYyOJDDPz3bEluH4F8GEylOILiFFkeFBSIWpwuVw3hWuNgeNEI1Pvuqy3mL
HS4TQmb55Q0YhCgcjXNNGtQctg9XWOMUe1A/zVCZh7W+necbVeISaQyGALuhlvu8kIaZmOPQmg6f
F70+ewdXJ4m/XjjcrJ/gLOso6AMctLRu1Hy+q3ez/OH0zyP8iMsCxg97lLHYiyTr4CqZxOfx6zPR
PuxUs1o1N2BN8uNgyaU/wa+RwS3LLllLYXLdCTQuEJQU0vy5K3gzcS5/AIs9Xmj5aYAlZMNxbkYs
GtSLiHuoop3y9Go89qiYPA9TMQa8zvRLAGDVsK7fUFzTAj8HK5/JDar1lyN5mBUijLUnlYctDscR
zklf090s/KByjJN1RUTILWyn+GLnzuRs37UuQLXyvn0q/xbP3llqetdm1mJCqXHp/7T7dF1moDC9
12kCvR1GNt6q2R3w6dfQv4cw3dMOMwAe+403re8lyiRnEqnLcgLkmKKV5gya5nWsBaNZYCh+W5Q2
Ah1CukbivPYBJvW+zDBpbdg+GFoV7J9vx1hSpLQdlOgECuZaeUhmiztZdoj3lEGdHhpyTPiuAt+Q
nhZerVvZcFzAz19mv8aCQQ4glMpLYp5MLSz1Med95eo3pTzlUgljkS8mWTMueaSno84L1hy2TVlX
xn1IEcR0la5eUwVGoGEThRX+6a8vHYXDO9wFRjPxcHUO+B1Gp/oODfkQRthS1NtkkpndQzqIOEqF
FtqeSf0QvRYW7DZtcs4aMYv5Grx6HCBuh0rg3Y8XhPBPHwdldfVYGgTV3QP8LbeAX3Y1EOJ2oi2T
oJpHctOrvW460DMzM91hGOTqTj0dKWa6NE90ef42vlujFzB2e/XLbDDIL2Mry2myG0W5OCYSGcqp
N4EhsM16nfuGQZ6irdlHGNfV9YyU6fF9bM+qzVJt9kGrt9sQMAJO/7ZjiTNzhELHxNIfqFRgX5Ni
vXdeadq1Ld+a+4cj/PIqus1BIjqsYxsJib4oUkvhtWfx1yitPFiKXWbP2RZ91N0Lkyjag07RNWD+
+WbyoYd6qACABfzgz4XH5EuyurHNmjHF5CVG3zISZbB+YXk1B1evvNgXZrIwkgrbiU7RtYDqCkzy
gJ0rtyiXy3yEx9K/kQx7k9LQzc4s8UtSq3Fyu3cckINoEZdmiA4QoWYVGkjSFJPUHynAqkxG616H
xZRg/n1ENmH15LUME6Xa9GrFxegIw3/aF7UBrnKGFgp56q61b8CNSCjTzfqWZl0vmC0IksG0L4WJ
DPXOTclF/JB0s9V49mK1DTm2YmZhhr+JOD6GoYfAZXnUeMy80Iv0QBB5gfBOxne+QC5SNSxaTaxM
mfuS5TenU1T0mogN6EePzZQb4y7jL5O3xI+mkZ3OQopqJrGauSH7aWV22PtHL4nShw8q6HVnM9lD
mRENf7c+YWxoTghLeXcQ7sv8KGgN//YYA71HHmmWtnp8HTOVRkClJ+QvsDZN1vLCjSdSIyvlbhMN
a1vXpzgesmWMt2nRB/KNNWzEM3cA4lDH6AIcIOhkcw3f1up5t7xzoqQBpPxZvE+vHDBtu5HDVwBT
M/0YKVdExw6G1fRVFDobiEO0Me/Ascd+X9B1qNtyZpb3E2LdDAB2w6x6RsaVwPlYDP1r8TEWQEBd
eQEUTDydKWoymDfygcLEEo1f5TP/mSr8Z6Z048YLgNn7vvGkpUPBH+ZbsheKdvFbBQGtT87Fgcsk
T5RoNRcmLZsMiPlWbKo8wuZuzAgdKanOum6d+XBh/tSY2wsSz94cx3QnGQHIxycimgk4FhtOPKNW
+hcFtxlNFV0XwGkUpv0i8/2mSQ0cpl7p1ZD6LicgNKhQrN4Pu4ai7dM0Zpm+1Kp9WccB9RKfMHRL
V1BrSgXUia9drPEihf6l619Vljeew29/P31E8CpOzAmDwlLsI6NoYLk2jPA5h3OYXW40sprrYHSi
SBSwkOcURSR/B6vh2Dzb3hKhRvOvswajIievkSHthkRStOcocy3HHxLDaZ6O2Qj1+w01XED0eBPZ
54xogg7Z0aclpp15cubKJXxeO5OO5PNu4plXNLvA5FmSKEiL35icwowPBjZy9Qk5wRSoRY6jmYgu
6jLUJdn0g7VUrG1cU3mLuisLyQb2W4Z1CzzlNTkOTtqIDlVy+woS+BkB17nTkFbC5jb452PWvJe+
saeVnp/I6BpYu6GrorFgWpGq1KIaIxpCaqf8O/lyIfdg4TMdCGfQvT4rWOlkiV+5Dcn1OQxUX3A9
Yr2ndGEZer1pQbr0alWUZBvJ1Z6BWJIkG67MNJPDoWpHLtl2VgvdsUG5r84LrYPWPglgjw5V0qDB
41DU/1YTA11bmGwIKkVcX/2zRtz1NCCSaXAiAImQi2jV2kSC7SpjLwzYMVCnerYJei1m/xj6Vyda
rcKuQrMlNbNW31pvzyUcE9NpD+vegidMfR5I6Kk4zQQUHE1p2tq+Xqqq4HLqBKw8I8rAoQ/4HtFD
d21lftNsMyW568pObR+5mggR4tzUXvlQAxRO2ZqnMtKU+xPZXkN4VKqPtNxzz89kM/KGqw+vMPAi
snyp5RBJp9hRV55zFQMSX4sEmmbUPJLBo+w3OQerq8ppgINj0GH+JrtHm679NsZ5ZlSxhjdLzFts
EbhwksPNM96TdVviHq5vkO0lksafiL/NiBomUFT6o5v5y+QHyj2yCBrdQEWhC8+CPDaaQqX166k4
y6YQFpkXV/Y5MyjHvIH4agKIM+wmXAvpkK9SsqNBLqbqUcLjX5bsxBW79ON0IxmcIHq4pJeW2u5y
FAWYZKwcBwzNT6IvhDoDKEF+N73cGB3YcVP8MNF6wlIpK9pyWrK1EPr1uMJFig2Vj3NqApqP74Q1
BXSWuPVOUdj+zB5MBShL6KGHnogYXTO0Shz3Ux0StRlj7osM61WCSR2yyLXo01sXt8cAwn+nit78
C6maaHzm1PHpRlkaG0drLKRv6AdPgtaYNZsfXZfYml2YHv05+FqaJoJz0+cel33glpL97FkjzhJK
YdYvBwVAs+Arq1udIyszOdWOpGi5vGqdgpg4kQh76E5+iFbbXvx3x/H8ZGXa/dnkMGXRPRe8lAut
JV4ejij8JMnwpjgJNajXWjoawilyn6m46u5SrU+IkMnBjMSmSqloe/tYzUz8aZAApKtVB2bJKpyL
lOmHUNGHtjHp3L/LdHoeiulYYlqr+Aq9OZvCrIdE9xe93oFRgvjn2n2EmPh+YPN7y2siRdSPjCXX
sQb6F2B1i8sPkVPR9KeelbSzmBrAYz0RjGPhTeU7tO7yM6igNjqGkTlV/32n8j9GBxBmDzVvvCEF
QGwpuHD+qRWwXOXH6ZuigLdvgaW6FKxDwM1GNJIF92zleZXZiPSv0PCs/NRXXbITGHq2BX5Nb9ti
2w7/7Hh6PMTreQahOR4X6DgpJSZ1TM5RZ3O8pC+LZCNzXz3raNLK9NW6p/qS0F4J4BOX9gWfGB2T
Cd0e37+HhE/0Fa0bN3gritekRvQ5lJVbLkCf6zYNK7oTvbzMuyNmExX7NGLyIfdtbrfxxbMwmKwS
YpyGSEAqar9H/J4w7XqiRhJy2FWhKoNRMIyA1NOaEseyaVCfMG1n77aV2KSvThOzf6j+hHwLcjOg
/xNZzCQh1zXymxS3+AhxjcJwliJWAU2lTl4lMm93gpdXYrhvDZrofmqCbUFtO92YC5v4jDD66Ssb
Lz0JDp/dT4ahI8+ie5toDv1UnxzOx0XmkBDZEv3RVVc643l7nJAdVTCkXxP32K8sGCmTMSykO/AN
k6pE4ungjvAnT4cvAS0cYlgrmP1wCD7PTuH+OENFNbpSpwOkm/KF1NQ3uXMQqDyW+ENk5LYEtOwF
cJcOerogH71yJ7ELGpOZ+dEaniEJrMLRNNMqkZfMqUXCirwYYZmAiTztWbZzfvw29TVzWW2eevd6
Dyz27GJpBDTvsd1cMrJP1rDFyleOfPRfR1Gx+kZ0Nn/MpHKZ5f+DghnQBFMFdQY9t82wlK0T/uwT
42O9vPGKpRpWM2kpCkPnYgKyOFmG7gq6ANAh7M452nDgMQYy7IU7QN5lHKjhCj947Nnh5lN4v8Ou
Uglgy4n0UcCdk5r0SiZ0UPPidIU9n1js5gtKTKVkCIJRcScG6u8iMU8nl2FM3d2vyvx4r7kwN28T
qEUE6MfkDTVyTal+3RtSZNWl/NydPqYv4b6IwLcrvJsdVigeLFqAh8iokrvYwh2zOFNHRQhq7b42
JrxxZ9DBQ5gMMgFQLtXK9Iv8vJYa8ota9T08k+MRl2Os5fsnUzP7epN458KRhIhme1oyS8kDSE+w
3yLNNf9xZ6FSF+MVBPLkY6DH+RRBpwDky7NtqNvOvP4J3P1xjr56S2cZy7kZjKAr2JbkAUtWaF46
CDil+ROoFaBqzLtHrETDqiWBaVwb9NJ0GF6oohUQH/vnJW8YIxgfUqV4IBO+RW4ALKuBPYw2ocmC
eV7lJMDBDXDVH+vgXawbuD+U3T47+Xm2IRFqeeGB6wg/7v+5KSdl/+mkN/7meq0RamvGcB4CrdIi
s4xtDM3cdBm/W7eaF+lp+nPIDfF+xBSstmjzu2RzEB7pS/tD160RA1bXLef4cyGuIbnRihg7Cq9T
fKNBsuwIPH6DtHSwRZx8/LA5Mkv5CZowaX0KylrRnnhuj88Dh7FK9dXSaZSc3ZVPs0ld1LIOF11X
BXZqPGZM+PjCfSs4sIGpJxo04nlUzOTjAZ++uUnWmoy2Lx/EHK+T0VgdWi/2gr7ebOHLjBiMXxUM
ZcsRKPt9BX4TZ3jzZ3Bz/AT5+ECKgWAJcVT5ZONFZAtOZFoQLOww3n9UVaJmB2GJy4Gaj7RIIBIP
I9LJuWPgW29RApzkDjhd5b2wxII439fn9rO99HCPtXqJm9ZZIC4CAAP95fbVoB5JP2lbQtvg4h/1
WmhoU4xx85VgM28qXA/W71SQMI3z7irUvMVk0MmG7ugscd9KEdIUQRAfq0FGyKXWOWNMslu/iQ77
NtzFplx3pd9ldqmFDwNWRldQG7wa4zgjRjLkCay4N/EdnpGu2GHJwjTuVzoUpZCJN47zmqPrPsxX
a5i39Q1U6NVCX90BHBQnks2vpfAnFOelDf6cxWgzKk7iB3wymQz3Fj1McUklhgcr3tMwOf418LB6
m6et5FRKspen6PIh8CJNa4g2Dw7iwrIN3HgwKH596eWHaKUIH8SztZsCNAxVWakPa0U0YCbO4aPK
nY3QveqtuTj1I6w84Z6SQ73dxTTzJO0DMUsA6ve/KHqpFyptHjzw/4hhplzMX1GB8W7B+6rjqaqy
epVUj06ADl+aVqz9Zk7ghcCRMcj7dPHeEZXj0A5gjRjNLhtVmHAJjN4/LeXimKguNn2tDs2p/r7g
IyttQstxSBiBNST83Jpmh0n5J7/+qK/zd8In/DEQza0G1yGJIMSfkUxtCXzpCi75yzwtmF4HG5Dd
G0/TcdMFL516pXs3+7g17j3BWZSrEYahnMhfmryQJ8eUqzpMfOOa/C2JfAFuGdFFhmDQRqDk9a7g
FsKYNk609IOkYeyW14v+oztfkdotwCRWg6n9DHZT2lkKxvneatiLtHXBpleOsiB22mzcTa2BuAhC
b6VYLMDx25SPSbpbvphYBY3OTIqobF7PKlJRkbNql8wa5ByJe/EKW4CDm2HJg+3k4OyHdGgrNsJ4
CQq1zPc6HIjvnx2I9RsOmxCsvr6i7J2ua06RCvy7xmF9GpN68uW9Smlf0YP7a2f8wVgUnvDh/7Ap
wyTGiVwQejzHkutczKgqnFyD28d2nkM2DH3ieJPZM2hWX/MSM4qKAfdHx3HMQrwA3sCxGnN3TfII
g6a4yerlkgUE5MKxN0OH6WikTDt5sMn2quDYa1d20iMGulh7z8wxfiAOYEHNcwvI/ds8tXQcsA5J
oYpDzDKGEpbFOfcxWyS2Y92o0lIFpyv/dGpYhNVSQqPGOIVzlfWocSOQCKU6tnVnMSQl3JyRA54L
EisT4gjznZQMeMQsM4cUtEN4/39/VgXTn7/rqjmrOfY5ZBtAOFVEzMPeAxdvi+5YTZ7J9xTmaRVT
QqXzS6rpWbSjp2qpMnsm5hyTRKIMeyvx7wDLXFrTelHFWlRlUVwSrq05ZuR2IUd7gfYD7msTg/w2
VFFv7xbS1sHYOltWzLfEtRsDYjFayBwsCe8LEcvS1u76T2zTeyOIG5DH3NzD8dCVECuf07aGXPSR
2tVHfSpFl7GJbLhx/+y+IkrZw9bUYAqjRomHcaq8yzWi/ecHXymY/r8kBGgKFqms3T2I6P7tfen3
uYytz+F118Qfd2b5BVoc3QY/4JYY/EFD1i3Kwlw4/itp4so4rpmLvLRRyEga36o8racng5kJAOXJ
diD3ZuG3rHV1hZUSLoh0Io8kd3LiYYyor2VApt7auohqNEma/VFBq0mpK81Xtcs7QC35GdpfyAR1
ekg2oZYJXstSB/MA2mAro8sF9PpRtAJ/qsrjmklZb7zEfMACrC30eYHNwgeUYJZEuvPQGjl37hGr
YQP/S0/DcVxVNRG22PgqpD9GvCALownK7qbsnoV5SfHTzqBUI/hQ348WoMr8B6M9ZCULV874CnSL
KPnRoOU6XAots42FnxA8iJ+YABQVCFAbFumMKvE1u/xXrtzuR73Jk1Yq/3D7fTlecKPrOKoBJ+Ga
gMkCSIBi1rEiFgoRE4zLi8OIKRV2cynHMV0y3WuG+qsgewQFP+2GMGZ+uis4bnPgpImOJ8UVO6HP
F90EKoFuRE9HaCpOgJXbtI1CxzevCQEN811GFB0avONzJppJCIfLFGdLO7moPoXLgrehADsXu27i
w28xSkquKrIkAHTi0HGznu8fHqNoYM5mSwq9XYiJyzoG04WmPWWvQZkdQfytnqg91W+yp0HSuGUu
R7ChZpTglu2/mSdmwM6Agaz54VR8Bm7cToyfDP4lCzeJCvl5ySo43xvkr1cjk8XPoViwiOCMEv9V
D79EF41fR/TojddxCNSL45ZMLi/631eLRV0ZAuKu0IpfVwsJDRdbJ21xH01c5/Aoc2NruSDck951
5rVet07QfeVakUP+BJnFuogGNxvTkIv1Mm6ARoWfFHYJAfaVd14mfpQaG8QxSTMrNaQ8Pz96N34U
6Qufe0PbrJBlOO+HoiWWm4xlSipQO5uDhChBvT97K1prK0qI/q19cMEimiLqmUq99X+GKrNGIrg+
eE/7v9WEbEdZauioyA2L5H13D5pUcCxjTTv6ZrAZP2/38SvKhS4ME/V/IIIYarcMFX4ggcqSyH4G
5KqlBOpM1OsUM/KR0cvUPNEnaUocQKL9yjjGfzAbh63+eZsSE65SVheddsC/LSlGsItr/MacH9U8
N6ttAYJjeD8xluLsQAKFE03OBLX0CBZe8DA0P+lOnVFh6TAOSzNOP9KVfzzy35QjkAzisxh2kDAp
JHmw0xIsuSLjMSC7JYnI/CPyfvbwQAY/JStWVRK/GuXFozht8vFpcmWSTGw5GNPRLpJyHeQnDyLN
KNmqsklqocqguVsIWNNztKa3rdUrFD8EnRPdkYRWdYitpYiaCknBzvIgXUvE3zn4jEMESUyV/GM7
j6EYhRKSGKy/LfFa+YYk6bP2IUsScZBEt7E1+Op74xwwotGe4RmR2nycebQKzXziDKHc8hSjcQUI
paJ5ktOV8I92GZ378iMUozii1LJWf83cRYR8u5XQ/qT7gU7Vtn3U9pAdx0zqTale/X0f4wZQo4V/
AOHflF3TZTsPVX2jFZFewYm30ZYIcl3lnmXHPhc8wXEUIbuwDmsPb6AoRvL1cl5GMbyw9ffAbkv5
3mOuWVjqyUWBp2hHjleto+GblXR2+q2ADDN44e7LJAwOrb9qYPc/rrGjJJfsCO0PcIqJ1WFRVBLm
dgJLRILiYbNz2lRgVybbm88jl3gwMFmP+gVV1kPsjhDuoskMz/B2TSUeu5ilbNSLQiQXP82jCEa7
LBO9ImF27FExjkEuzcpdDwescZYzQZOyr98wksQYStyXC22ZnLZqr45edDenaS65WRlYKVlSimkx
hRRijrlN/pASVqOu1mhVOuhFH5MOxpopc2wwyptC2RIvEdj8bRugdAuV+d2sv8cruYuCw0xfuSkt
cOpYEXm3Y1Ikb9mNNlbTn5ouChvdH2Q8hl4l2z11FHQNQvCJaafbl+O4Dkmx7SftH6nl5Z3qrbeT
2s83Mr8aatfNAPQu5QFjmzWdOf6qouFUY1+8q7jVKZKp3aCziN9nAnvuaEqSe+Pz+79gn9km+ZuL
pbdrmTT+ZtMIbSNxxlmcmh5a+xdNbm9KojYpyoYCcQTngSL39IStIoy8VGuOlgdywzngWbdTZ1KU
dR5euAr43y/Zdkzr87A0KgwYagvF2KD87+CFDdJwoAEWWf22xu+0CwftU8TKWZjPDjoUzg/UWHIa
FbCxuoObUBdcvkpvv+63bYK5ejapq/nI0WpLSCvt190xWPGJZhN/uypGePL7Pavb8bZDAZvBO41x
PWiSTXf8k7ozICiNjSPyzWA07CsoEmSMhTybDJ1hjvLmdux/rE9mAXFGjN7rSSUOPwISZOCem+N8
mh0mTB3BmS2qQ9tnUYKivHc95ZZujAejgOUXWHyCi5d0lm/vxLu7hGhWQDN5NyvRU7DOld7nIOqw
hMcdbZkgXnlWhM5U/OcYEEeChOASkQ3NZG5tfPPLWLyBWoZs5SPMVHiOFKKIk3Q9zxkuygDYn0fB
NdFRoNaxw5E6l7RveI9Q7IHE9t1H4IIkc7QxkNcRE9bUCRzKBRuKOEACg017OoH7vUOZy85POCj3
4uPagfdOiKoR0bi5uYfOBzvJvrrmulEaBYKVY41C//GcbLyULzW7exNkywzNxno8Cs9rAtFKRgqq
kr8bQUlZX1KhAkv7z9ABf/rhwAGEWQMLelwVnMCewvf2jdjjYuQ7kiiRpGDydiSMJnCtkS41dAEC
LSQgB1looUIdwSroCon5rRzu5AD7Kdn7FrqXOxPJa04FxbHUxTvyWwnspwdx0Wc6iWldV5IcXOeZ
KjE3Tt+LOFu20069+JS5ZfWpgmRzE/ijeD+gShTA83JkA2fNCr9G2nhYPSx1PRfEkikTjZMwJ/zk
SJd1O7NGa+kJ136VWMuS1QomJz0cbAjlTxYyGavF+mnVFdXCKzmasdA7xlXcy5ICo/tb29HWosWW
RTqjuUmpRkC4CiTrI2kStTpzTFtPnyan4e1B+3ygahV+/O9Y4n1qBNMVhC8jlFq7XW5HaS7sc8PT
ZTxUOA0pi25Yh2QSivP0AbrLsPaE7SUCCFrEeTq7u3Gm7kzCg/BgdXtfXS/Rw4Z/+gfmbtY2caNa
6gBGdo727EDGTL4FgusTLuZ6ipgwSI6Hiz+PtiWrCeA6HjyrEh5Gdi2ep+LwVRaCsl1gRKznwcyS
Zowp5P/WwnvZ+XlgCoyahlc80oHFShouhU0FCIa1gcsgRGxCt9lWbAod5GNmVk1yImuuScrjwCDl
/asmIiz+JLVmRVkbjiAkAxDKEhbMcmW0KbA4HNdReQZp4zDLWYKu9r66/QPzwAyHe+FSdayDzR3X
Q9nvnnqDSy/ADY3P0Sizs+WD5tPU96Bj8+xg42ULitdaJGCC3n1m30NayS9XXnc6mZHvn533Re+w
qavbQIXT1ma+GzioFjRSN9aPMGsRwD7UzYXzOLMCBMVEbIubueh24sHbBYTIHuooS3h8Ss8NVPRQ
LdnP1XQmpeVXXbNgojR2xW3jZL7YgkG1OdT0gb+3c47od5r7aABzzSfYBntpuNo95eY6A9CzgDoX
Huh/k7qFU2QS2KPgeY1T1gdsm+pTU2aCkhQ1OrWFve9i2UX2zahQ8dStqEFaPMopJz/thvCx5u69
BI3ExKZ0hnxMFBCtvwo5P45JyB2DlSWg2gGWYOv3/F38z2YLvyuqfLCD+lzBmIhjTfEQglfC/ean
QcTcZKjjv2jQrNywF9CMSn7Xms9BDkuxxKvtWwEMH7Er71+Ct75c2K0/Ekt7UGsefWCvrz/IavPm
omKbwc5Yr28kfF6n0LsiCoiEQieG7FA9LmOa9trcd9D/Hnh+hPRihOqD3MUX69U4DAq96DXlsXrA
AM/6o5J5okD475XwjZxBKyFxct/RijgboBi/n4zRhgJMW8dNQF/4y7KZRkW62cLKo+lMZUSxXFFr
+2ndVeGYRxjYl/DVBSPouRppyJqcvAOwU82+f0neU0+FePZu2K/6s1mREWySJgjYdYDdgOJg3BOr
0WF0qB2lPSqF0QnBTq2OAyrc7l1mGm9pPohSKqlEQSUwOvgpHEh0MjudOmV8Sz5Z446PdwvnMLtc
3gewGpeAXntaWw1QKhqk1sa80rd4aOaYEQmPDrmFFOS/ShbXMNBKc22VuoYzDxG+3hdnXiSR0pXQ
MQMsTkv2Irhf8PyVMAIIQgLH1WZz6i805Vl0DeVb30oWTZXnOaT8Ae6qAKhDPWrlP/X+kv3581ZE
yMhyfrudwTH7TcG+WoJOH9T4oi/VeU5AmZTfCkz5GVVnBO1S9LZXTpkwws0TaeHKNY7WiFrjjaDR
HUiY6RrO7cBuRwyWUcWD9P6AUgVz9ESZlzFC2iG5gwOytUTr14LQhhQonPaj4mKdZiAkBuVznjMe
QvuR7+pQQl5YEo0K/Zgegs9iKamrDsuVNrQa0UWmwL8ZGGndwuD6iYI2pB6HHoWv0JIWuB9hEDeW
5LYNzqa+/2e2RzYWVoGyqNml2H1/wu+RkC7hD+kYiKtQRCjW13TMpLqbYkeLAac/jjx0vM/1gQwU
oaQHUVJy1kmueC/qMMAneahskrAHI8nfXsaHKzBFfMG+gPZG2xP8F/Jp7FVHIffcRCsoi1LKvnE/
0Ow1+1QXOWMEY8q8YM7dLdVdqCuXkuD0Vt9dG6Ij0+5USuU4DpmNM0xabV4RZfC296QC5lbiEwyz
hX/355xEPxf4HsS1ojg8l4g2VyQ1il6ixkpKlRGb3G6fnXJ8xdG93pNphFkbyCGQXF2KdpCVljF3
CkcH+gmF6mwHXtSArNnv0fujbaYrdGnKx2yeK28RGXuMQoumGhWqnJ1GWyhM0TR+fNTxfLOdcyId
vD/4ERLaNrSH9mtGvlgf3zbWwJwhU+E6qXB3FPqG3fP623Rr5S2Ew2F1Tj9Ygxz1XLDeanT5hHKy
2WfiDdWiAzI6NHfRq32j7keLEC01d0sMlCVUiTHJ3v9Vw69dxaEAYGgxBUpsYfrWuMGJQPG5WFOY
5pgvsgKDHqTewT6tl01fE8aKYBM7rO6DvR2XUzAbo6NusIRvcf/TtFQNxynk/hrHi+3b6wMz5Tm9
iSI8WgFW5A7BpOOz8mx+msDB6osX8pjMTKr4/+lpiNmqMDTpB5Z+McefvfyRGqqgFjvEFu4ERA6l
esO3yQQmmdpCDLvstAUyBJhHtHgn8h5Uk1sY7Qk6r61blfmgnrXMSTqjPRE0dOmJ5UpF9abzrO7p
UU9kVtxxMFwrbABZBImn398hdropz1Gw05gSYLBCZyr8O/8NQ4oHkXjxHdkbWDwmsOsn9CKfS99u
+SjPg3tQwo7kfh2MziZg5iRbZISxvcoHf6dy2p6tHMG//AIaT1kpsnsMVfvHyvCyZixXPQVZIG+j
tD5SbZp+ti8yq6ZvQrpy0ALWynlsUnL7Q6gZlOjg6ZLud/8UIFahbNh80EWwUOAUIH4LMop3oLY8
61A+xaCG2YRcj5UUFecTzjFNUlRBxly7mINfU9DZtH8weYO6qzJ0pWS/719kz/eVKmRWkxFf7vB5
1ZZRcIbVjfqh79ZzQEifCW0eLo99FbyCvJMDYLnI2eBklWvsMtmsaabTiDFD3SEuDB9nJ/SUyFmX
SVphKD3pMeFg83dpi95LMOmISfvUf7inksj1LHKGQh4Q0b853Ccov/Mu5B20rHYVHdjECl4ZAbGa
n4M23yg6oG+wRwSSam6ouSP3/b9siCZkSQXS/XDv0tnvuyGuf5PAYBHrUQBhe77G86kyWYHolw8I
Jmp8iDIcA7WuqjJ4fmai8h0S+DnGoFu0nLL5YYIBRTM2oXpeISdlEgMyuDlACDEhhDRMMVmT/Wzj
CjRRzzUiy1u96l2Wt6pYwy551yM/L7RKS6AAnv7JcA8uhaefdv5xoJcfHe+Bm5jvbaA6XlxPYwGN
h5u1gZWhO1hJUOQD8bgXyMREzWfDZSnINVNW3V204Yut1FNf9gQlY2q0J7R8S6XLhf+pomYrD2BI
4eHmuT5qOBkDe2K5+FjujX3cfS9wCe21K6YH3O1IcNOKMYE2+FMchW1PYa9l2Nug2Ulyxb22Kyj1
YsZdkE6KkX9tKziMbdMkTVpacisF33Tbn2JBVnrejAIPigN9I8FqVdQdR43urkqUpJ+mdTKa8rd0
rWCON/rU6iGEETWv987JQZ1rx0Bj5Esbv2Rl6AI7CpJljHipYoh+HVI3Lb1XH5MGVUcFghqYQhrr
s74UvbV2r61bQ9+EtiI/zu5O4iAjDWkhos8qotSvXO4eUAYqJR3sJGtrnnTdjppkxFJFw9vv8hfm
KEgfyZ6fBgcwmjo6zE2P8YzFy6daZLTyMo7I+rkV7lJHX7SM+WBR94h++bX0+Yf/y2PoItfEu43Y
OCr0OHQ3Cany0vEMyWkTp1b6AsP3cR965uI3v1QR/04nyGEWhGu7oxWrgvefncJdLI5mhe8xeoxG
yWRTdORt5ZV6MULU93GCIuz6n0dzmP938tBIwHv6cA4Sx+1vT9128UFKjnw02COgY74Uk/ITYeG0
r7RSVNTEp6UZgAypR2hrlrWjlxxPQyJ3qJMRx7vmL4Dv0tgKRik21i8P/gLv9bBSycVjviy4yzUo
7Dr26KntHoQDSjbv2luBe00DtyYHr+Pg4EfXcxekYBpS28bEv+rJ/t3oGVF9Ww64Sb1KlK9cd5Sq
8n6ism0KLcEl1Revc7seadvLALOBitPgErlpRAksdkIWslNSZqz9G5XDRxC2bf2fnuk+N+bMNJZQ
NV6hqCV7hRQpdXCS+XMbc4AKKnjjd/k/6i2Hd+yN6qfctcGhS5J4ioADVyqA+jpH+u7YzaCEl13g
A5+DKx3JJwlFkDyrP1gx+5ec2od/cNDsJmOmP/4F6rLRDpC+bzc27evCYzsIpxrvO2WGZwfMN+nN
sKs2GUGerB3JtETwTvUVoshStBBdk0lckduD+IHQkLUIZ7ONs2H9HjFLQxX7XpZ9QKjp09qWm1F4
FvSDXi1OUuOIQp5qXqYco2YAJtkk+WDZ8fkdYdIopn+9N86kwf97O8o9WXrbklFqyIxqVqhSxKgz
Sn/ckYTITGEMfKkMTtY0evMwWN3ftFJPvOvovkKfvX0FO3IfaPGiVmgKPmdw/eclGBMwTu6T6Lqe
mgK30BHjWrGb4kHp9mA0fzp+O88MMnPDI7p5nTTmnGUqLp76EAItW+ssGkpTd6Kvygsa6refvx/w
ItUwqbmRV+gLBlB26XhyYmgb+yYCGQaHPwR6NOz3sAcC1P5L+xG9RiEFdJsM94tT2OsCMQ9KyCcR
BQv1KOJPuWnDq4Om6dEqW5aGl5GWkuwtGp7a+v4mhLTUC0c1c+wCPTEUQi5UJuJS0G0lTE1H8B6N
izhF/Jxcu7XdIigXHWmwFvHtisSPaAE7MPMoOdfQckl0czH1akW8NGIZcX03YXZHbvsAAZgvghjw
OoIz1C0pWIhR/XKL1N/Est8UU0KV1JoiouqyjjDVGN7ktSiztF5IT87uDQ217AXqsaBamw/4WhpS
m2rI5EDVKimd4GcxM1nVKpV+iq+wvO60aMTzPBzP9pIEs8yVRJ6kGsxLrrZ+S6b3owj9NGisvEZ9
t0lVWOkr4QkI41ykDXaH7w8uVV/BWW5ulGUlLeuqjkCQgRK/H2FyBeuy8MHMDSG4I/j9RNiD/ceG
Rk+VzqnLX0iZhY6pjUN+pFQfnh6CjSYSS+SoI6UMrFr9X8zuG0jMLSGziXlf49VVxfxsdMUDuIw5
/t+NvYShwhgs3tbYPf/cMjrupCyQIcfTFNTUz2xyQYI1SoA7RJP1vSgLS+T3rxMfeztcIFYS0jjK
WWSi1cKIZbmcaDxu1PM7jQ5771XbTwCs6wR9B+0jlx6VdAI7Ka6ambpsQOlzf2JJCMjWIgyF6BLb
5ZQHHQ052xMxcfHioQ5F4D7GmoGvNiX8yeBmMPkY1OxwIqtsdMNoBQEjLzsmW7Am4H4Zx70tijsY
oCCRVis/YRIpRBQ39dxC0joUZCvAedcj7rZELQDiO4NhkgfkTnJWnxXusgXJiU5GNM5Me3xBc4iZ
4D9Z11h3CZIwg34nrj4Y/htITXga6GDbljK8kFIK4fZqem6suUGA/UJIfsiLDRasaWuf3W8gfwbZ
R79nz1fQkyIGJUOPNVCLDJmZpgUrr2Lq+23f7SfDM8kD5jhJpFD4yjHQTinvFEOkD+chzmPXIIY3
nkRS0Wdbz3aODZLZJe2bGjJVcKF1qlpQxJhT2p/Atod8x1jvt1syoZkWaFIw/Ps+KoDbxfgJqo4N
6djuAclxD9RttFaQuMi+eIzHNZr/1EKu6cRyxI+DraYjjIfn7AIgJ1HNKy2Fi0Mfsrt3R0bL4x+i
yiivj1roDuD4C726GYsQdw6d4WGmfZEbz4crYTcjk9zBWRMOQJfA4Hiw7PGDGZbFzoza75u7LTaH
CPFm9RrJGQbMeXWdhH/T29BF544p8YYfxRFmSlswIoz9ih0oS+FggCzkYOjJMg70gwFRxq9ZUfSq
+yTyi9wFQ46tkzWB4CnnBxYwGHVTJb65ineeUfDL1XF2dcBQJe+oRz53ddQrWz1JMUjqJJI754uu
ErfBHe4rG16WKXW2rnN6sUQgq3RoZFhpbzUpAxMI7jjtbByvab5ZPg+VXkU334eujegpNQsGOAY/
Px+jUycd34kF+CztzXqiAjQfxRAcUx0fnDkdsRLKbnLYvQg4QhOC8VsHBo/mqqSIVTpCcOIUJeMT
V+q+Nk4697DS1zIc3OSI1QFdvS/oFcU7aqPAsV4ZnJDFr7EIwntwVU4/3ERivk68b0+PxV2wruAl
fJF+/UAGfGf7EJfnWO7uSDV5bEX7sbCVa8bayXIhNAFmnDr+NrQYzj2lZ4UxpOLAlL403LwVOR50
MFY15yQn7Tb0EmOcimHYk2XjCkv+lyQXJd2c1zQjYJwldfPYpL047+i2bQAaQ1JzT7979agyUlZV
ySuxfXAdx4LeQ/kyqlyD+GWNmB6Gh15mvhR/oR8tnX8MlLtkrCCfDVQgSWRcXGYqfJioMcLK1hwW
hhtw+EhauzQAtb9manA9oBQ1QJ44v28xuHs2kOU0hiND1Ob91KtHmtESV2BP9rtdT+iV0AunZlJn
aVPfsLOnUEbyG35htbpILR6at7GPKI8zRa5kfvdMQ/wSPukCG1I1J4h38pjuQRCATuUtlDJaXb0G
VU1jrG1m2h8L94jtJ1L34pGIA2eIrgI6fPp38FvRNxhMNRR07N4reg20mxn7jPFR1V30p/dGMXuc
HJazB12dwxzgHkvszR2gKL0xIA7U4p1+9+7TjbYfM1gaQrbONPi+HXZ9XZRdkZaLwRhpw2g7Tr6p
1WRxs8GKp2yuOol0b4rGcl7Nmh5EsF47F0ruxKMPIeASLJ5XF6p3X2jmCicWU1yK1xu/vxQQ3j4r
xjlgRwH2R7SxK2CKMyv4FK2oiVEwGT7tHyQhMIGHBFqY48Oz1Eex8Tv73foWjos3Nf8Zkj/J+uOG
Ei+4IJEciUmuQ3UamvB/mCGxnwXWmv6IvWdaRwWoAeXyclLTFcMHYSf6dCBq3Z9YegPq/iQ6bE0w
+eIuRpTdT1VdkrYuvWNeMmj79L/QHQFCeloMlt44JCo6t+Tauo5aHEuUzr3gVCkqe/cO/AnTyq6f
HyeHwkloKGT40Z4jiks23q2IB+BzdltJr6BDn3AtAKRSZxa3vQF2CKyjKff/fqPDs2mz+ma8L8U1
KfMuM6fiax1AjAiQMzJ0M10ejBj+wz/WAwn838vwnUyTgRqCF0A9UdBCayrZxTJQVhbFM5JYCxga
nc3zeq3sNTQjarcX3p7ImGIgu7biyHCtYbsDf6RK0OdoTFWZrriTyzQJ88LTirNCDxdyFjNSItjq
x69ew7sf0q38a0qv1d5mxaoAngICNCk/Q+g2blysqMW6FzDisE7snd+rHFZbe/84dfXEJf/DNfQb
uRqCtYRPZK5Xx/KTI6CAYq1fhC8aAD4Mnzz+vQTenQECcpDJjEIJ9Tav/mOhE9uQyrfIeH4u9LZL
I8nStJwti5a9CANLS4QVyNHWFCttQ/P6wjvzx2w9tXMYu6ZMnZ18WHwElahvoT97IT9JucSqTHZl
YidE10for6mO8Hd57GQoXthHNhTCliMUaneHAvU4cpEdZLbgJHI/I+En2BfkvTDguQve3HgFFq7W
DUeGwMPzCliKC/ggEIPuDF6UqVJy9LI7ifYYIEnXH9kESbbIKRJo2gi4XnzQ4Z8MOrwFinlrNcK8
yCWkxO0nDr30uhte3PRxhsgZwZUurtm+KnQblyLpmHVk4azX2zcB4vOwKKRQ2IaCAu3bW/xOy9I3
AkuOaKq0G5IxNxk8upTp1jnGc0Ji8ad7+OwP7Qgifcy6LgUkvLp5OCeHX0QADZZymo9GGoCpyiFG
te5yR33i382QCbiv1HQqr6/XLWoyYEqUTEGoI98kRsB2RQx7sDah1V3IsXDKxvvH8pYblgHQMWzq
v5W/vQkhqC7xbTHoW3BevFmOb4VgHj/R6L0h4HlN1lTgzLqsyQDkqkkCdRzeJFV600+THGLLHzbS
OVC8Fn6MYzaRlxtjK46kF6WAIA8hz0RMZ3IV6iYAvC0mJyIJs53KP8paEdyJsZXz3brDUM7e1Inv
rJEGPfVarRCknqIgq7cDVIe9hq5R5Ol6qR1Zl+jAj1VR85ySsGhD099kg0iSuFvXkmEDSY4BpIZC
kdjOBU4iltTrHo20vX425bpL+BRar89MZIHzm4DPB/vj/H4XUxIm3IAUID4Gdl25DGPqu6/Ou/S1
iD2F55Xyx7KsPB4nJCm6MtuE18hjR2y/SNg5LD4exZLH/5M+dFLWa10F9Eldh64cnu8hy7uhCdc4
ABFwn6evZUPObFkuCdUSPEJ3BeOff56eigqUpU2od0d8Aysu6JlM/HQPbAWVr96ureWCvIHn8njI
fAFn8Gz5tkfwp/aZ4Rbk4TleXMtNd7ACTJwHQ/ekebZdWYzP2MfAq0NGgdXo2IDSGGIJqRzh/+j0
9OanTIV6Ag0gLhcMZbfTNOUH2KClBEPTP+K0EIhZI6k7oWa3HN5JgjpHkZGPc/sFe8A2VXBv0D+v
oAlfebzkpyigIKHWIXIcQ+nuYe07EmrNYAQNQ8iipOY90zlWRk0+ZmGoynrnVyoMDLkDTMga6bqt
zDEQYQGEOiANUQhjPncLU7B7fIVHlr1QbFaha+7dQ427H69Rvc2ZVh+rPVzMgEf9+OE7FnWOjuH4
vW5wWWbgRUk4th+zowPer3B/IPSu1jPu46nFJVvoPoxFiSxePThvxropaZMfoZE9QkH15sbyXgb0
pMaL136zkeNvdxhZUUYiVa5eaoMhhMvqSKhJao/psw5VdQG/z+penYj/DCTwdlnEzKzCQpNbNetz
2frA3HOprkivEOzPPd1VKFatNga+mq+lqH0Csgcck6b/goiSJJickf1+99fwncI+skNfhlqwl7MT
SSksTYT24//2b8pS6Ufq+oCx+Qm81Wvg3WqZw0qEYrOvwV1xzbCJNa+16GPO13jg2YDRozcMolt7
QCiJn5UH3LX2rWRY7MkJWbKpEXz8vfyNI0G0IpfVj6e67J5VyBhshUOogCHR2EwrGTfbRMKHg36V
rw+kVGbjm1vVO9SODpokeFreCCJH8sNBiOrLLmZbBvZ9YOOvF1zDSjb71LEvDHpnOocjFd92OS22
bZWZNNZGHFlwY7uyu1XbnV1OkC9ldcEPdWTlccacXllJw98jAcNx/HzMxJPDQ3D/ge2MYqHMqql6
uDTYlMSebI1HAbF6fGLX45VAtMCO4TMq4YwAmIjHGwRqRxfQnTpd6aYS08wOJroJOCIpXvxskul5
1uVq7TF5KLndrEAgRZTj4B0rIBC9iAztygUMb1BPoXu363R+sA7gsykAEJRICUq2Fg8mFc85qLsg
B9sWfy7T0jgASumeuYttEXS+ADOBM2eyU9o9n3yL0CpKV+RsvCFD7x1/lmc9nE5Qe6V3JXFxcNjp
OStvunFbUZ8xdeA1mQdIQqA0irqEhVxUPz/EFkYaAM6WYCXgBj1nr2XB4izUmiA8/A+C2Bixafg1
tTVY0hi7xH3c6Ij3l5dQW09vDgk4uiw2YMubLeSnolTB0fNrZg+IvRrjJEgtFlz2qbUmlQqi40u2
uP9jtlv7ojRkgSHNUzXP3jjMggNEIgxVq7KqAaeNn+oS0u4K152G4cZfKUEmEUq9/aynAjaBaovw
8jBhy/AVslL2xkULHAeLxf2/zLPZg6L5iKmNMmT0Ei60Zy1BFG3qa70g0noGDX0ypsl9UEeRitW/
DvteldeabciUgcM9GKWpGIUXbjmYsF5yPDeLxs6hOT9gkBQQi559Ro4y++/c3VvOHQeSTN0x7iQk
T/HBhL+AyNfmZsCN9mBSZbGlFDlAh39YnpBMSU6F/6rq0EAx9/kv/wZkuh0AWcun3hXdXmpI3Kuy
kixnkXnPAB2tKXBbAdavBtGndkJCX/ttYj2TNI/oZ7AEkxkRy5dZY/mjGw2dpzMuJCbLSEzb1RAb
hz2/X9799HwTehrP+1J0W8dqtjaxnwhVWRaZYjHVvBnUvkprkOXIP3wkfcwcQV24c3JJx7nDkIY5
fQ7hPrTeQEHM5Tcg4NQpvPgp4iNC8V5JjsGS3qaFIWEK/MBKNlWlpnRz+jRA0cV5WdEo/g8OvDI2
FSka9dk5ihVC9ef35e+xIBFLOPWucxOnftI12Q/s0ZWe73rMxqiOdDsZ07gMrG7JXHU/OZytYNAV
jRYE5gGI62ud/REeCWCpGqN/v110YTfXLyEpR3EVs/6VGpJUJKQqlb7HpIQ7NnJXPEemJOHgYGgf
dmjONtfPAMuX1Hk5npdYA3kox+dsjVjG9N5g/2GOQgUYE+3f0Q8QpTPpU87qIJr1axJ+3+7jfSqP
5ghEm7nTV0igXLBaZy5+k7d2aDLCywnhifjo0LizrkaZmFzU2t6r9MqFOEPPmtepkKnkeHatiX76
bKiTZ7x83ZMc1TQYBgjKYbERO2cRjqqC3MvqjymYV29xYHJRBYD3uZMz45OBoPLCFBvN92XU1oOe
Xm0xNAbwh5pymq9vmImfK0J5Q4rRsQNUCYnECSqE3KgTGJg2lbQstlzJYZKz4lPSe7xUdCze+afJ
87/nN0BMCSQKnCA6dfYJDAFuuPD34HQpf+TIIM4aLkm25ywh2lvkdgb+7G2nClbbDt/Al8Q6u4dB
MBW5N0UPrqlIEYhqyUwZA7IGa1bZQkl/PVcw89/Iq/k78JU8vrKZoHBvkdqiAvOGUykB4HXW0qF1
bgq5Kaco1viR7vGOv81gaP+lJCw65fLWckFxTypQa9O6fcKnI97GNXyx78VgDYH16MVsOPtc220r
D/ckol9JiDjGKlmb8c7IFVNrD+6REsiiTxtkmdXx2wg1MNy67vdAS5QB2gtpaezqmfem9eKYRLl8
F4TOHoGkh08Xb9x/9vutBts16N7bGKmCSlgTO+ABK/NJRSbWceRShbbWL4VVOWyCU4lVw6PwYG7Q
YiDeHF0lnCh+j4/A+K5fLYmMiVKH2oXCxoKhyH24N2JS5AeNS1eMmzIDfXukiJfGKUuQxK6o7U7w
yhEv6f2fPzm/euo+N4fqdLb92e7EvSqE0vrP8uKj0427Q8Z7Il67++6ncd/tndYEsQWC9nA3HYec
1kUMKi6rXLFrjivyVKXMKYoCegXQHyOwem7dzTcDyC5pB4FaqbB3SRrcesg/yFahMeTpJ4IspYLN
CKHcej6EUc09rfkocLjEUDdCExF81rx543hFVni/eTR629u7wlwyhrlGuocgJML31OImpEIdU9GJ
JQWUcNpYDH145bB5jFlE0997cjO3A2x1zI9EQiPFs+cl10BfLgZtYzbXtb1yiBa1ZYuIrpEGSU05
/AAlhjgYYvVf9Qq4iGtgWsFmAVgzptDrPq4Yp+4vm9eempTDOKD3Vr+8Syq4c/qqRh+8rZc/ufDu
y2qa135q5WSeGwNBOt36+jc+0HzZ5MdHJflIYxNYp3I8eLlEeBD6sdNirDXTNiMqvS7ngmEi9cNb
zT2lbPw5M4w5nT6MfefkG1ixDGZFFyN2zI/xjoi4Pbk+FnkGplQJUgb7ZKtAbFm+LTyc1FfV8FjF
6aFawItOSUcOTQfwCJ7aUtFIgStpiiHIYveLwfv8WdDPsJcs3GJsaoOWbG8fGRrqDh4AYcsvzq+j
QizdHVqmQCtbKnGSKB5pqm3mHrkQfFlXJQWO++an5wlNPj4zZ93ptU+ZYVOHue9cAZ7+DrH5b+Ak
mzjCTMvNbYMTft4sHtQCvJuNauztFHjhGsT9BriggdX/svc1y5PCXtrrcgehIO/6c2rIXXWrv1t6
XzvnVcHmW+/2IQphoa9XasGdiqPFzYtDg26PlEJ24i26BM0+w7rs4nRu10VYFh34lpLCKxv1/LWM
ulKtDeJIQ4HWqihRPpo0ya1IN13xD+kePUQ34+MiYzz9Oq6it0WeqbUBLb2aIcYW9eyMOLv4oUKA
JlbTETgior/bND5Ga9HF5AITWzwU0GLNAW7bcTYiuXG95X1rIu2nsMLatzTYpm7GWQNLu4t7rOnl
CwtQqWGs/FCgiXxS2Ff5nsh8fMP16b+Ep1xpv15Y5Y/lWAEXZ+i3nMZJ0PbnLrAMghpoEwOeab0J
d0t4CRVNp26soQ208LO5d4GxZxgggMPqGxNFQVjJYTSZiZ1WALs6RnKXp06oVmnrB9J55VuEnGuA
MMHf/as/KAOGqn9Y4xMivpc/AJUE8YomeTzlhyfjJP6X2U/alyM0ATHtK95UjBrQMZP6EViLQdTQ
q/yQqaMnTyUMKM/25+/Ika7eqr5dFvlzO29T1E0aSyeAWapGc4Kw5ASTzmzEKkSXz8J/tBO59vlR
jgU9XROdcs6va+N6xe2rYhj2irKABqVK8LzA9W0GQwBDlcKd60PA8ZQTsIXw2eJBGWNV7c6dbmlA
LYB13DoJRjaLoInU5h2Ks7sm7/hvKVhzkFrAVeo6f8HFCYHJJAm46Qdo7bfsfQMnmyORS9ldyX8F
NSA2IqLDtR9k6HDmwucBWsBmL7dbibwHbyZ+ZRDqN4phIHVdBF9ymWNe2/5A8EI50zWMqM+Mhv6N
lwBWIXcNyIh8z/6n7/zmVHOMEGWbPucQhjuBkpXtl+cHd2NIcW2pBAQSKDJtEMVp5bBZ9rH4U3Ne
fiShSjwFo1vI4mlKu5XlNUJn3U8kgGGmYrAADZR2vEImVXXy89ZiI94JVt3HGQBP9lSfrdxN2B3S
cFkd6aT6zFQHY00J1Y78Q9B45j4Q+FDph4Zy62LCMnS738FaTBdjVNz9/D9IVBf84CK7tNqTMcrw
iMxEOw4cEDCQMuAtawqTsCVVyPCaYz6K+m9QSSveZWBec+4BPvGwvhQ9WQ02SYwi0olaQwSL1luf
6qPGWS42RV/wTROKwEamy7j0OA1m3nArbGA8d68RlVX0hsSi4ghuL7rH2AZ3tjMUSeWR1TIRXuwV
EOkOcIHdfSUXpXp/7WRdTOUIjGMxHR99QKJTK5NSuuCdMDvtZ33U7ff6tO28kpx+MeDqi6bysBfh
gc7SMvmRqldRE7rzpwEtyD1qouQSTuHgYEGeE7eLUFEpKB+uZRoFY31U6oPJA08yEyvShhSqhQh2
DD0JSgM0kpYNj8qAbg7LMXuf2NqLe0fcjsIIkFNCb874UWtGEp4v9VuyrgTpl47KMkdEFTU6tRye
LGKcNvooYyh4ZLBByUvW8Nllbt2ZFh2pA78cmojZLWnZlLQPdosPOad3rPucx7Tiiev6RSGNlUWy
uDGvdkFym0E/shBwVGBsKwhkO8mI0LEhLwrgh94LZtpq/QlLfb5X0RKmE7QtbAGtPb0iLihcOC8L
4Rq0GYP9sr6xs0mJSuT61u5X4tvFqfHD8qQxYHq8DPNRRAErAuydq/diiJs3FOAGbHXnHdEpD7FY
lJlJp81Zcq1rmPhb/G7tTfu7WpWwfXFicSSUISV0rCvoHxwP/EwX05kKmIpNfcgGcLtmyR+F4VL+
2PHI0F8Z2g2WRl98BlZ15VfTW6c253EuIFt2InR+NsBh7AVpibMVvi+w+JTbqRlNNRTkVhjdEwUM
pgFHeTYDUcDwS5/LJLSH6YDpe7xqvXdzlGrcQTcjBx+EE2dB3ilO+w5Q1/ScLyeB6wwVfjQHGmJ6
C5JIf0DrxNIbv/kVL5pe/nG0C2TZ70M7LFVYBepc/B37LgkaXu/W9S4jt3DlN/XHubYolLjc5Ren
UJO1d58tRulcRxRu6VFbVyG5bbRjAuJEkFNLklsKSZ9hY6xaYfFLmsCI9e4+fPAqnKM8yURbPUvA
PDLd9xOdx24QkVk7Ehu8vp14U/P82y1n926Q9enDGawGU/9bAOFu7XH2L/5ck20mj4gqhiIDCWyT
nnJmN641bZ5cO05rLhbGI1B/IRQvM9tQrqcQSGC+8wW2ksHKzb566bvrePIo1RlfFEd1JJlu+/BN
o1pt2AIAjKehw5x0lE72JDE/LV5j7ExmLEzFewX5E0wtwSruonCP3E9FEENHnI/Pm2PDCmohbQo/
WbqHHxo3a6tz0U/jKeNVd99XxOg2g2TpJz2Jj80gFAht7hViTzsS9RDBFBqGAInBs4+q7hT3EGqm
YN/Nn67wYh8KC5bXmZRBPokWdemgoZaFRRw1/9v6UPT8tygIzie9ptxdZQMTxT8MNJt4QQoXSSwo
+UD0GThZa+p0t9men2YiORIMeOUDzuyQBXwyYxJb8g5Zl4WpEMB4qmfsGlDnHRHOm3o13C2aQMV9
e2GZ/KivNRHjtFvErKMI6/Hkiikc6xkXT1n+9Tsv9jhGrBGC9Ph4v3e0V9dv1yGH13foxbsYItjT
TbZsKUCZ4UaW9WnLLjMosvWBVmuBKOW6k35/EYr8HIQWjs00dJQU7aK7gkX3eRmQ6nyMCh8XEvXh
rgJtsx/ZILMz8UmlfT8VrjhANBovp0vt2ujDK8x9WCBNrgnQLF8A2QUa9bWTwewj5/VcwAbxPrq0
NBDSb3mFStp+WGrM+gN1R8Bi+KVrxMgkdZUvHafFO7oKrVwH+EFcWnArNr7004N5X8wZQoKTFkpK
/DkDr6XZ9b4Eni/0pzwRvu4ZQlHuHdfdFQbIfbIMu7mw9LN1e8U8vFwWIoF9E7mNd+PKegpKKbfO
xM8EUuSI8nHrtFeCSZ3Cj/0SvY0Ts2c08GDgoy8Ml6o8m/ZPYOGCD7i4kBGqHTZD8ekHzUFw9y1s
DYARiW9b3vhSHUi09KxxW8Umi29ZzQXNGlqa78l1TXQeleMxBa3Y4q92ap3AR9s2S6xS/v8DL9UE
klr5o4Xt0OVD/9EFYZbSyFpWx4erF+5udxuADWn4jW5xg0cl/HJDMEBvWxCPi2jq75GkTYWy26Zi
wrb69zyB5xhpcsILxDZdgFey1h8+YYj9rys+TkjWSbFM9y6rau2MRokGskjfLVa+8kb5jLrPxnAz
bySip3wVRV8uD+1TVC6aGiJb6lMm0sz9SDesWGRlDPjWrH94rw6k7yUUD6A8erBGE9LXNzvP/PJQ
7U+ER/Rv36LN7/hh+Xk48fwfYHQZVdawKOZj1MpXxZi7+UifG9rnrvZqJWbU2tnXPtusbs2rJG8G
hAkD3tNfvR6w1J/joZgLSMTT+Dfahflgjx6Y4G0dIQUA2XwmP9qdNacVLMLGWLJK89jD2c+T2SDU
idEBF+mbzCAs9wY52I9DlQPM4mOOYYm/elpd5CZpi3RLBwIL8UpckBMjemS2YOmIZKL2an5XAMkt
XU6zJjRFLudsyaSGbJk93oa7D4wIIHVl5SQ9nPnFRu2v2jECQvIjZXeNKnRHzfakCGEoQdXo+It6
fbNMQRU+sMcLojgrToZ9IOgUdvmhpETZGLUPRuMZivjxsN0Bsx8JPUDZTv2sriwK2eInaIhjLSCN
fHDE0GuKusA1I356w7W3NGN+qAbLIRivEiC8jP/zJDbDvuI2/skMVqw6SzLlq+fF6pZTJP6PZCj0
GoT4p1Bq9IboFgKdSioZWTeNQTkx2wJCZ9bzexU2/q9NCK9NsNBq0xmwhJPyhnQVWY3rMfL8Aqim
VghPRvEkBrYSn/YuayLgnxix7BnTBmbVAsQYJMkO/i56Ck252rN+zB9Ao9uwmFanKo7qhYVBbgI1
rK9/JnicW+6LUNH5/WAKSKA2EqVAkItNqaNnlZ6yOHSdQBEYgup0jZ3GGEBtdhBgeNo3DFWZH5XL
Y9Ffcl0foSF4xE7HUtm6j0k+Lr0W5Zz6shGfKO72ZyYIlhGZqNdFT3BZf/7y/AMk62ZZIlB3iJtz
dSOUscwUwhmAEMafkfQ4fokQGNP2ZFwutfTe8g/P13DpYyGwJFjg3gTGluExgXVMQ51u8PEqu2tT
+sUrljlcgFItXUNHaaE76x1vCJvywXbwDXe86IfxMqzhJeCpWS1Cqqqr5Il1MbV5AO4jyxkaM/RN
wybJFYbURKrNz/ryU0Xge8Pdemzqam1fSmr1OVhi9bgaYdEian+x63uvN69RLTQyBj6XHdTZS5Ws
M4qNFRUIEkULS8wP85sWc6CcCIKeC0cUmeCrg25pqey4tiNr60jZoCoVi1ugewrV/h1ewjdVaDPd
2mCAN0b6z1m92c0xO8+tYg/B3YSsduIbAGDpyzZdNdAy+al2DqMDm4DGDCDWSLf78XEJBxo5xfqP
pgcSbYTKuj1jJO3zIcOQBmClydnckxDZCiFPp4MiTpyqws/+36cq0WwWzUwj04fE8h2CZuCW+iG2
2qgrtE24EbvAX0/h4/rYkDlqHrPAnn9lr6ihqFi2+2vk1+XNz1XWahN21z8Uq3P3VOJPr3AFvE2b
eu/d8BjpVhL6baC99la3HXkqQoQcg9C8xrcRi5ZCpYdwq8sEn38a7IxfKH5DgItbA1Y03ohR8D8y
DjEklG1xfi2gdxCkAkOnXklLKoJ6k0r0gIHcJpQ15oEYt0NqJc4w3BDp/5Oze/SSAMk2S4qd0dVs
iKlG4HuPV3hYm/5KU+y/S0fPYGSTL81EZcp3vam1SqpE3NkqNwzyq2l9k2yS7rYSJN1xB/IFFn/I
yNfDauROErE5Hto8S+UudZAuYYq1JdAF6sWf0GsYltJVIa94m8hZFwizymP8d3ucA2fcbEzs6jD4
lr0EsIcgvky+p1zCW6RjVTjxfTrEXavYBS6l48rlTp82FjiCckxy/3HbEJJ38yh+rRSUWioX6yVe
TBFB6WANydekk32C10PAHJWaQnFczwg/28/ZytNUV9XKFUgvTpDIneUTeKOgPH07tKktQQRH14w1
vuDWF5KQ3Mb4NQq4Wb/n5/c/keXbVpmVTjV6/GGeOwuGiVv9WO/eaV49N46RR960Yeq99XSaHZYS
sXkrhzhhky/QHg/zTXwZQlcliKpTDI7rrxPLo4w3Qy62lD+B6heuPKVVfue9EagsWiaMpE3N8Mkp
k6CW5NSLaO/B46e9zRP4ISXtVgjeb+b0k4Ydl47mhcfb6gF9fJAstSbef4qOuqP6b6bVBGNPt2fm
8XWF2jjBbHg6UJdMsPfILK2iV3P7ZnTtXsLFC9sCxNgeNuJs9mQdeR2naqkfBUHX8Mw2RpjIxrlk
SygdMPqaktUjpgOahRzCHT4Z/W8obM9UDfoAZnRx9X8ae3ZAiVq0k37r7Anry+2k7Ugy9EZ1Cjz5
kt4fJLABnZIYmppiplM26Q7mnqfEC/oil4iQgp4NcZ+a4QAcuZ/XUdufa3lXYnp461wxOj5X0SL7
cobSbcazW+yjtfD6nox3qvJdX4Y13s8Cp0Atpzfdq4R/ORdUVGw93K7ZrLPw9l5mcYg4iXmyX/jM
vbG492x5g37rLUUIkrG0LE0MaDYxEXRoQ81LZaerbfbWZAD98qOUvWHwDx3EB9hId06QULnbyUV7
veJv0lKfXC/4O16V8J4xw59oN2Rw2GtIRYhk7nabOlvV+18nUxjRN9QocAGe/7QTdlFgv+90SKSV
N73qll+Pc+M4/LzfD0qVDSlEKk2ZHPcC1w7TGQCeXuUXjjKTG2blI6zXW/JFhtblk7tz6M568c+W
P/zpSzH4WFPVIIX++rnkfP2LjrT7i0I5pFYLW0/Pg4uv1R00zmNvY+TaYhVJySO1nYbUpZ9Ac17K
6LAxQj9lae9vaytNI3VBWXKSX9o1HAPr5n06vkylMm7NTpELVW7nJMAYe19gztEgJCoft5zClbSY
/MEWJ1u3QbiAaJZ7R7a8/4ibjdCR0VIA2iBqrUFsnpMKP+f8i1NL7UPBo8IfELQfKFx9ArG4BQI/
EqmGwCrNbvs7/5K3DYbOf5ZVgGUkFmseK1yqGjr+7QDkgb4I0yQSkfej/pfRWVVa+GMnwapNyfe8
4xCEEHYwx1GNRw+uMZMRdB2Nuf+dv1PUYu+9Xo4eLqsZEMtuNzbJXv8vXAlh8xcQ1STOyqYn7J2e
ghNrrRauoM3LPnENu3aqvHP4UePY7RJxmGTeIocYuGCc4rG38gANYEaJgq0Hiu4o8gv24MltXRAC
mQqT6bea31AHbB7ULEBIdbUkobnC5oUN21ajtxnFmlhw74Nsb9Uqpcvqfmgja5La9OPr2Y/4MKgH
ez1QgHQ+0z4ialBq6IGCVXl+10S5Nm9JAhgXH/Hnl32pZxkqDA46dztJ9HqDo1MNNnxjfKzMujRg
tuqmpoX+kLIHv+OlRj1ZNlnX/NG55nBn1xefhdgTBs5GzQ+cZGhHF0GfhIIEtMvJfZoP3lOLLi32
pSkANV3v9FYFxcVf9c+Ax8pce/p4ZIQkM8SrUJj8tsga1L6PrmO2+dCyb96Jlojqqvhxop97ETyk
yKbPZUJ4MMyDXBwmuUUOIp6ppR5h/oD1Lqu30S0KFtvawVjasd9TXpXuVF9QrWSjGKQbuT9uejW5
wZb0g9LlSmdK4XStWiSOS1rcSmzUDwevMOT2ry8Tihy4oD0vla7pZDMzYeJQdPFyDbcUrAiPY97f
2JiakXVHd5T6gv+n6zNAFEfkUDcj0qblbDVNteoRSXTPq9b1lrdMn87Ql+am2tQDLwK7dyvKd1va
8zr8WSf7QkSI3k5st46pcJWaj6smuAWmn2XiZulBAandL/QyUWPP4bddz79dYt9EmyDgn73zLUqb
6a5IuqFTY8VrCYhMZ9JsKk0hcwc/xOGXQrJE9mkYbtRA+A9c2Dc2sclY6wxMSgtuRYK1ZRdBkHOo
JlzjmXN7GRT4jzJRmZhqpw4VlGRSheF7EawZbARVPBzkSU4zWdLRurldCwde+cp1nvbhqJVeW14s
p8Jkx13flJRanZ6dzHwlM8B8i21bCcpdM5QFq4om3Auq7OGrF995VsrCWrAuoj319mAtHyBKPziC
BdVtpPBGiK+ptAsrnqVPwKQ/v2znNbkBf7CLbjeBByK9WVL4NFxRB/vEBL07lBdyuP+RoDeNcnkn
c+KAqC25fMhozY999abphdU0KWu9/ahQNqSZyYSNwCrulKne2f5YeT0Dpulax84j2rn0ScL1c1oz
+un3+fKF+KTBgAeSjoP58j5AGP8MQFIYhtlSnNOokAH3hLaAj2svRgUxiJNPQuD0P12MslCZmrfc
iuwqxV1UnNTSHS51G/7wzViHFfGzwJPIN85XW9+FfdLG5mPBjRo3H0T83AVksX2w2Rta9BXCsvaC
g7qRMwBPdZLv06ueY4CdvADwfAuUi0BeLipkDqBDcE/XTzgqvLTXvNae2wYqxq90VFBLHOdi74vB
kXj+raI2O2yFYTaZ439mfnbQTyvt6R5fWtcjLuMCpqD+HWg/8Qfq1Lx8slqMIK4GLoisbYrY3xbP
RYqEjiNWNAFfULVyeT+NC7DVKeg1U6K7J/ui4viSJd5bW3q2oaNrR/R37o1GY7FI6yobfG9Nq10u
mHrhV8ApynrysLv7vPkJ4gfLUhmPiCXIME+kzVufx/rHM3wAh2QZ8SMrbBHF4Qx/VTzLD33asZkf
17Xe+CHlRBEAd7klkintlEmolIDPt/gQYvfxMDxiA1Xu4gkVYUQSzwvWChDNAjZDkuHXmSqIUTPR
LIkxIvGCaFHuhqeoR6O0orduic3Cza9Nr+SvmVrKAlbZaWOIa6rBVRa43NCuXqyW7dE5OlA5KsDm
xYy48PK2gveMcbw4cUnG7LOOv1E0VEjTNEEq0KdTyklxNgjVlUtveg+O1iEKrAGaK0/BMdk20s1B
QJtZqv34+jVq99z/jgodMHu2dNhrQdqqFGDKKgQgadvu9xhkhLpFoo3slRAiT2aSyD27iWYYugtk
iJgP25r75O5mVp5YHFRkV7u+oUwsVJU5jxRZqjRxTK+XJjzPomcJZx6tmCpi6eN5r1MmzbahuQd/
ktZW1xAyhSawTYYIbxZkym7Hw6Rh2LaKqbEFsujNpm1Cd5Ki8cPaoFOPjPD5ON6Mv9w9RRCZv/X/
bDQQMfF7ptzf7kT40V/eazqVDSbEPpacpBqJpTwsX3Ik7arCTvWMa+SBDIV1HWpyzaUW33mPW+37
Rtvolc3gRMpkIv5YSFmykIrUfCVTWSVHwHnX9stN3FZXR0+9rwfv5FRqXfgUEugSUgyruaStbr4R
ZnmXjifaLECCgbxbDq5qXEOlHezUdFkLFKrrk1L0fwHdIk5rryWtH32HNCSOw4THxbYgvbA5t3jX
gnCLrNsuLqLedUgGrjcY2pkQa4dr4LPhCa9qs4WUSt6x2upi+35MI2o3YylLkwEiC0jD61ggJDDa
+V+yKXKPqIul3pK1UWtobMgk6KORdV2jKKx/Y3SvUILpI1G98I1egQSVY0GGX1isqvcQufC+cNjF
2sPTx2ELeEK3/Yz1upYFDF23nqW8tcGGti2S3snO8KHBrkqxILg8v6Yt0M76oyFCe+KjunCZFoJ6
raNRqS0KJmBTF+5l1LrOM+ipBiz/ISqE6mgyBjMa17A0n0g8pwSKcZooDfQy+NdKzPyKIPpkhaUo
TUZdTwZJ1e/HzlWTILMtSZ0sqDI8CxqnELMGRxP4zCzWWDG6drCnwIDRKn6/QhA22NLzP0+fXDmC
PJblyuJk9DMhDKpSCOxuD0NfM2LU3/QtxX8TV0pYGMXynhP+susjdzqT959pMZr2HERdxfpSVTI/
XV8zsooewEXZbz9uPTWZ8FeCT2voDt/u4qsebexYLF8ddqvhZvd7p/23bNKChfOyrB9tehvBAZAp
ZVGdcmFpL2y5dMv8fDIrbQbTEZf5Dbe4l0Cn1k/Icd6A27nanYqOf9vRqJdBSbEnYZBDrFp77Lyh
sTkQFusX13YNGoZANSiGx8UkI51po9rcVL8gP2IAQXpHW2CQ72VfH7UZQddqiPnkEGaHhgn88CWN
fuorwmSBkBPS5NHnSjy1Y/o3f/kI/4KptWatoqVUXsK3k93BqTIdQJU9Fld4aHYpUdcoah79b8Ec
MnLAG+CywMu9swhiZDmHZGL9PY5a0jIMgAOXxAdqkW4sTlt8JzFXeH1nsXPqDtJYjGoXvmdw/9kt
oF59L6cR5IWkMum7GcOfmKJkCpMT45dB1g3r40iSJBEofGLQTSDn5wTdh5uUWNayIHALQ5HdZz/4
NVi73v5uXkcfoLHokp6HYva3EQn+dScI9VN6EkpB/AIc2UQeteLOplUokWEsKsEplLk4Wtu9rzR8
n6y9tzmvsWQOfuBo4jQVOgh4/U06I+a3Ox21ugX01vevEbesFHghC4YrqoGKtU1n0AFlBGRVcHyd
+kRfU/Lt8CkfIRD2CY00XcN6AMIDGHlM/+U6vAuFT3IfsqGSMM+owM0YaEzv3jnf/kuZkDyX20lO
KywvvV0PTG++624LlZNnQ5mNDOyHAxp9Z5LRCLBGU4n2S6ouxByIhU05C066EX5Hf2EH6F1SqjKI
W/ypmhuginBGxJ1mRCUhaQaEVimeyGFwbAdD1+EtjTQHX+0lFWvRgqQjUEP/ScZPtBWFv5akmyH2
gZwcsCSvRBSqlJ270oFMnddSYg7YVOu6Ylrd3px5maJ0m4UOLyFAppN4mxfatuxlystPQbETmffz
Freigy3Ztcr8ATqlB2EacyIakAmm4Su6SxV8ThU8jVM4yYdzy7/W68Uj7i+6DnI1U72k4ACaGaBR
gF4Mig21BTXzCGeYvzjk5TjIdQMqCWauR3dUh2OdGFSIy1uzQEXTEHOrr3i2j58vfIn2UvBXGqsT
6j17yxYzL2GjlyQaerzIYuXqr58cLoFOZ60kE1Adu1WnXaq3yWo5zM13EiUUEexXmoY2V2WX6vxu
vg9EIq6KgNMXbampRxTSX8W7PJt6PxjZyQf+PHs6GEAYdkSnGmCQRAFerMB1Q0Kezome8/Czfsh/
dNgrg6XqLIMCz6P4gfb1uGMSLl7sHqh5n1xWC+t0Nj4IRRVSzVxy8dqDAJCgaomTK5HqOgtw/vHQ
BV5QxpHAaT6EFR7a0h5iDZ0q+B/mAdHZLpCmFv9w6K54yAxSgvgYDTwbcsZHLSKK8s4mdKq4pk4w
z+YiFl1iJj+v3rpRB3zdnm+7mpDIcxh1DoL2xjNMtHyBjClrmRLR8MVvMd4k1sKs2Zh/fXuhuNDj
h+Q64WuJ5O7yFMFSI7xyKNKz9i4KDayFdAYUNaTmN3J7VkziRcVfmc/NBV0SsyDZcF2Gb+M/0tn+
qxx5ZGBr+y9eb7O/w5BzHdPvFnZdYnkxdq8tDRu9+bLoWAlEC0Ld/ZEPdvWo9qAbBzSFXUSBjq71
zFv6RWv2FRu7ifCrrokjYFvJRNnNxRcDJjOFu8JO+i+/HKBOtMVltaWhDsMdOBycUT59o8A7uK1u
nMX1yvUtLC3pyZDiuwyywFxKhY0xb/sY4nSC1qJ7i6YmuUjMiLwe13MO93SpMffNkxnzTM+E+/RO
yMHDJlLnPtWlnnvgiQs4YWTbk8ooYlWK1qRn8a9/gG/mpMVbjoXCCIPW8tHjIKdI+0nSkJqboUhE
WImV28SLV9uOjm2PN07hiwU/VRRec6qUla73ikaPO/LWS9mo4uctjib/CuYMOizmrlfEp/Sbgl4f
rxgnZode7vSvNRrcS+SLviLJTHgNjJcIBg59GYEkQCVtZghrnpTL3VywzdAv9w98+dGuOm901H4+
lyRaW3OpIYS3jkdi8TNCZnNVKW0wWhB2GMdDGxwDWItRqaFo3ah8wXJiSt+vgy9DLvRlcy8JSUQ+
jYN6b2A0JLfSFcIGkNVdCzpGgF4Sg/spoKFGor6+5zjRaQMSk3dM/We0u6nkajGh2108d/BA1IJb
JIMrtuJydh0IXW/Mx2YUIVYUZiEjnL2n2JjxIEc2CA3Y4beLQSc+6DSnk3M/nFKQ8MR8TFfgvXxh
W/BSyZ90Fsgom9TyK6GaLCbPQZqpoXZ51yHrYo44XTB3Rdb3+5hyEKzDzdqe2q3xs84Khci5hEdd
oiqIKZcpJwn8fKUGLk+PmV7AJGIy6a9rcrhQHrrebyVpNCmouxHldYComsvmd8VkgdPb3PXdTg5V
WRq5s97mJWKMIXvtDIfAeIBE1SoIINxOkU2zIot85T3+B5/iZ7b7x7WTqh1x3fV4jUuOtCPmGqZQ
lgUxEpwlBIssrCKwc2gsnV5jfri+HPj/2Br6S6zEjcqCyRBondIy9/2NYZIkev9NS/cvOnmPjUkg
kMD+jJMTs+QLeagpor1vGqw39F0hcHTGLUSByYFc7JMty8CnKhr5RWJFukGiFcJK5RWmACgWCCKb
bUq0jiWlRk6PYq668bISdtLrqv5/952uMfNSdZZ2mP1kOF6SpQaNHYdw81A5fhAGhzC36p5tU5QW
SCZ9vBv6yc7jgNdGY9pxchKWzlEzZkP0qZAyLPwc4/uRUCSJ2jD8DzHqlZBpCo0oS59j49BTwFLW
3GDvk/zsJYr2aPCutegXBlpQ43aWTudx8eO+hL8w/HiS1KbI+DfNRmKjJ99BFFA5zIfJJMQ+kL1V
tpQjO/gafKqr9Ku/ZgR2FhPGuPD1S64i0jik6lm1VcQyDLZEHPpjxz9Sk0AkbpcoBkfwBXxcBtNK
IDocuL9LxtKL3O/5hRK596na6EjPbTX6z6giHdRU4c17rc6kkWBRGnVMS4cyayFZabYkuMkvtKPO
bqa37cK8fqlflTKiO+5ySx8QwXtYHDZ2TLToJRQgAfdXSk3ZWxWtL+VgZO3poS8aiV3Ke8paRX/R
rr1kPMAzVmSSLUaexkoGmasw5cAqnB5s8oZB/pzRVUC74rq0K9FZESDxC2TNOkNXxJ28JKLpiPZF
jYs0Y8YwgBdkpuw0HNFgm7F01IqHYC1OuHnYbNFZUCbofgAFlcckE+L0vf+JYeNhh+xm619aGimy
TLasbarKRWl2gx5iUyN3vWdbgC2lF9+Hc+9/j4wE5NpFX/lHYIdUx0qeBpOZFeUF454qDsy2YDZs
D9p/e9+UzpqdyGRCsL6zwpLgzfsO1a29AwckckTFldsjrleNwMQxWObSTVpA0RwRE5GUb32a7xJs
UiCQ8N9MDBAlMLrm/DBOykVpP0GCfdpyadW+M+GHDWuSJzFFjYn16lE8RieXuCVzB8I/OoC80sFx
7+4WjcqRnX8qIRobl/e+e5St84f2SWicFrtOMrezmoMxpYBVJaw00tXogZNubEKgATtg+TFMJXdy
ehkShDKGyYcMB4bU+icNXc0XCqDfpRiDoL0DdkdGrBMHXdVrrKKvoldXnzi18E1Ud7v4PdZKDsre
kvqpExmY1MbXERGXso5gFecB0nYteEJMOEH21P8JKDJ0RV0gwdkdQfd4pVMg7U94pZ/QKaksnnZP
/b/UoFcTTQ6/Bv9Jx5N9wbuzQQ2ELOTlnW7hiKJFceGJc0kSz6W9X4twVJgXrUCQHfLvUeAV6FNp
5MW0REWQJctPZrA9DCBhLcEglO6Dhnq+Xw0zK4OeH2aoPBtk06T61Q8tWE99TWe3X2533Os6xEXa
lSfYm4URNt+zSCCRilNF7x6RopVFWqtAN0cz8CV+UowoIZ/Nc9i3NtDFWONrmzPyT6iUerKNU6zu
HCBH3iNbJKUoYtOFvFawLNQtdCn+5wG+/nWIuX8jS9xwz7cBM1pD1opG9LES+Uy5v+pz/CSGpfwh
9dy2dNKUtrKTziBGLt3ToLfjirW8NOjkr1FQIx3xEEAp5/0hKtsJn74Ci8lJyZU4QkRHt9PVbDJ6
/H9Gf2JGn8yEy1ZbYL+sXvxBthNjaVavtPRMk0W5SC+fyBlEgtPez2Tyzsx2JbwF1g41zLutD/4+
MVMM/y+r3EZMEttAwYN7tqlZU3rtit8Okrc8rKSkQvctOo3nsLiYwhILdTbKkCZhatQ4VAjxlc+7
PpiBmzL2DKMIdvkKxutd9qiKUfxdaDOsmT6xFcSl0doA0mWDsppZ4oKS0+ZEth8QCTLM+IkJ495O
J9aBOsOiQqta6qsUD1K/pZb6x6IWyW8Q58Qf5ErrQmVD1mAnavxiYX1/gHb/DOWPx4wWKPFmM/36
KSHgTutj11kRFhIuCfChvjNXCKaDEW5cY+SfLfVJ9NqyhT0PvhDfzNVH12LDnPq0sd8KJsJAQ9Wu
rqvWE8uinIzJ84ervQ9DkMlxHJqkU59I/quqAmtgsGefQ+T/AE14WBgCl9mCfeKRmEzchs3gutDF
otJ9rQ04CJSCaS9ihHQdveedX06ddss+PAsoG5IbWCkui+q1uTj4fINsu6Gs0JGFWrz5dAJo65Yy
z4zeZZfNesduVQdzrjAMPrB2V7RDfIUYl7pj4rL+CNCvtX+XTGaqrNXM9VBdGtDtKVyB1jdaylE7
5sbDjyCOuZBsRCVfnTjNhH4PM+geDbPK74F4O5MPk0wNYrCSmgE2KObHqUH2rponYpZKdLvr1xBx
5eKuRk0HHGpQAt9++uxe2wdb/oJm1D41MdR5IRtBF+0+d3+M+B6ibMZH1jbzzPYep45LUkwNWju1
Bj5BpSabMuIey3xq0K1cj9Y8FNc/WcYu92aG8TLZcDHLIqjD6cwTvme8ZiHoYxjrKN/+qyyNgEZ2
fmAkrofT0pZc6NyNQrw0GEN1U4VoL/QxmnojMrHt/1QKvOMA8MfcJ/zAgFQPT4Lb6iNQZng2jWBh
OMglKHgYuBHX6nCKivNz+kTO+EobtX7I9ABip7GsgGxmXJgDuviBsbWsysTGykFb0sVW51MDvI4E
aPvFAKRDQU/UAvt95smtICyNbD+/VzxmOhrvceaDdgMGumP1xOlG73N87pmsD3fPqW9goMuREo9P
JehUSx8EwqCOT793D6tOHjCdl2wpSSqcnsEZd4j12Z1ggUGa1I6Crxe5ed2He8IgTgzqr5gXp/52
/ZGtb5o6gomQvT/X4291bn8BrPeOOxqcK54vmuGtuv8+O47Uoja4bJe6DfOj3/nJ9+99zAFxEMiW
Zw5FzRSpPUk337amJcR6rnqtkw3rFfqmOCH8wQwzw3XG3jqa+RlzNUKkIZlkk47h4B45Cjenr0K7
F3TbjuILbN0FTT872m5UncQ7bKv6NIebSgkwnzrgZxv5NJh7f3GlK+/h0VhFU/lbF05wJoB87BzI
4HcROhdRetw1vYLUV1OEHpARuU+n+44FvgQuv7KBqOQLGxHpKTbNnXuycmq/JEa4yBJ63jYIVlmx
/1wFZX/EekQglwqVFyYFv5NXo7moDKs4m7yjISd2HPSsgg+lH2a1vY62q+RNi2aJJ3KzrENVTeJy
2KOYJeHzQ31OV1W8EhvUCAUNMKsM3r1pd2UZhS586wwKNlsOnH47S0uURpyjreTUC854JBmSK/nD
RLjQQHg4NIXTUY2PHBTSScnF8rhVZxAgHxJdyMo+w2k0nFKb2PF0c9QhZAlqT/zN0zYSF3NqqNcH
v8/GSK3id6FyOqNChR4nori3zNO6PutrLRcEUJvMv+2OteIsBBiveaKFOXQCrjyQP2RaHiFzXfFX
p96Nv/Zqby8WLtGZHAqBkoLCqgiBj7RvlCf/OYzDVBSNSdVHn5aWHRSgAMZNy8pUUeLW/ZkqYPKZ
RIoVsZO1tOlcgoH7kgo01jkw821F6vgvzQ+Ly26sqvsQLEbTvNo8EFLd212ZEu4u1clq0qz4bi3g
zppjxmQ5gs87opxXY2PrHFKjuDJfQnPjq32PznLws+8JyTZZsb+CsBqNZsyPrTZDpmxy5mcTvmFz
BkLq27UBdKe67/+40BykbkFl7lfhEs+xuOu4yatXqYPLt2ffiC9YgBQpJe6/takL2rHzsKUqEM2f
z8fqvuPGSS/2PYRWCloW0CFnAzNCCMR+aunWpXRp3OlOBZ40oP6NSwdfKKDAnfRLSlZlS5gXTQSN
Kg2hcZSnYqICLfLx8LBoCk6WbGUyNvuJDUwV/d7+HFUThlOLWsFC+W/A5Th0+J72912ck4cg1ZKY
uiZOHydtrc5dilArBiWzQRYfqPOLxky93953SnGxs29q4d+hpfcAQo5QqBDjHxfCtIA1FYNaPPJ7
KwduMy9mj4xdJO6++TNq2nq6OnPqWcPVTEUpDda/Hz4UGMAn5zyvgzoPfZA5mtpvKFB2+g4/btZN
U03aT94H7VJtjupqguPhIRhIjCQm8dyEUOssLScS+hooT68jvoitrjjuR3dVwcFW4d4C3eH7MMmK
HGR2X8SxJL7Yb7GkebJQHvw0mqaYpxptb4iZu8FOQ8WNzUFayU0fWz+FHGM/xJ/Iu+T2QcatSs/d
2QC88NHBXQzk8Ca4oQ1Ecruu4ICofFoKfKhYELdhWfrkZqZAY5jU0xVRaRPKP8siY7va5Xpcx63V
HMBBRCdlCvAjX09v1Jp+/nowyHYOmAhHLT+gpEyKUCW3Ib5X8NTS7dioxvFTpvRb53+DiDvET1jH
vYHA78ETw6cXl+gY2bLMIb9zc5gkjEhSlxnBne0sI2IozGz4+MoNAyVDr3cziUUt1dX9hlsA4FZE
dbx4bkb+JUDwwKcHjbFciUkQ/172ai9wv4/H5VRq0VmPaUU8DV6Leuuxk5vifa8WFqJnxwKK02QU
01yAcuJZDSeEgjkR2/N4JVCmUijRqeQ4JsyV8HWeURlIW1i/g5k/GZnsvPf5tIJmTr6ofIGQVD4Q
ir1/dfewxG1ul4bfWg8Lr6AliiCQZJOOxoQ63hVGExYxlmrDSpL47+CEqXtX3+IlUZ46re+7HDHe
LgBqVgpK2z0nkgaQcgV9D2x5FBESR/0gYOU7oIkDrLzreJ9U+Pp2D18bmnK5kYNfRRAxrawQRGE5
q/xoEEAOaxRRy1yGWHrRJElP32+OJ3lPwKajAhBF1SW8QdFcU0hvBW4HqHDsh+yYrSQAifbIIy9+
bmoYeebitiLHuy6Pfd2uE3B+uGuhEfYXl1Vp0RxMAX+yy0IeQHvnpg8GxBmEjsNeC9ouPts+sPBq
dqQ/1DPf9VxWX/V61Jb/8+gkOKisr9iyfMx+VdtaPvTZO6F83TApI4TIhPu90VJ10Ud51ItwJK1u
5IZZ+Cjp3KjV63U2aOoaHmU1Brfe+NESa/r4cJPgomEevspMl4SXkAx9+kK2SFO1nxuvQpfvQAfk
vP+5SB1McJETknHuRB61JNhT8CBrwQ3sFtV7CtDRxHjfcHK6HKYCX4/Akk74WXK10K6vAFq4fJiF
g8ndtxcam7b3eFNOpnGIA3CQj+E0GzlSQXwhwUZqisNvJOm+jD/nJTaIROhAeZgNXowK7pt+LaOx
d9l5tbNHVnxiQGnZhMO2DMKb+iIw0N7RxcmdJOU27TZGki2n/m1SG3WsnN1gLSYsoZ241rb/SEXq
PeQv5ufLYPyoqBZiGcpbeaUkQINi0rt6TwMRzf95Vq7xVaFCj1gM82eFOGVqcxN/ulTRs+8ahy2w
A1gzGQbHJviT1L3IJBjOD/mc5msokf+e7ErDSQY25kjDO4JgKOGVixqOj2MtDTlBViyUCFuW+isU
NYQGq2Bb4MZntEIX21iSFpzH8JSyYSdmBnTmpbehlFqiU/sQYTNmP78UjyQM0u0c0Xsn/tcrxDyJ
WslkUPoo+nrsmx62n1R4Y6FDSwkrbl5V0kHwIW9173dM8fMMCVPmcZvg19qhH3OcvBFsYMRZouHe
pgpwyC2wKVqs8/+VyP5dr28FxpmlfLhyVPmQlvRNqf9G+2MjSAGH1NMlq6fDMUahyqIFeqNTfJGY
kUUDtd2N+l2gaIGbGs6hiVjZzfBjoYi5O85oObhZdQOZODx9/EiZbGZnoGkVTTj3ktk0o3YPRnae
pNH4DsaVUA6E3QeIQbvRwU4kdIsIjwE2wM+JZTBpuDt7LwCpvXKFoXE49mpLXuzilV14plDhCFzw
VneKVwCgRtQWQx/WA8nwAZ1zbcbEWaHQn6YQOCynFvWZc6Y3vHcRgz3DgXwszka3HnUMpj58AJct
BaI0TOLdZWFDl8wG4MlEf7P4eeXYPIIGJ8a3wDXZlU7Vd5rBe0HtENlb3S/BsAltbAyPvFFMUAeZ
Q3uYrsjPTob49THvKUB0C10mneFIW/F37nHopgdo0mtw9D3nIodojbCoCCQF9Fh2F1s9p0zHZ2ib
7BuJE9DyrOeaud0EZ81rBGlHMhwq5gIVy5ZydpEAcyir17bG0kZ0Mr1+6X2LJuYYgzcpqThid5zT
yiRyNZDMCL3zh7r7G+sN2VWYDZj8R8ypGj19W8jF5eMhjubRtl6cmosUMkECVK8X7NFVQJcAZl51
CZ8JUuaZumBPEGfRKxnKumdmDchaKOGokLDTS9QSFm3mDYeuUWF2wPHs0Zae1pVuRaXoPpSe/PdK
n4Xm1sQP6jfnjhwGSwbYg+FZ2U/tConBCFspNARkuyrvwmVPieqVitCh8x5qzxx/4bhB/7f9Tmsb
Ez2DIAB0Z5OAl2hSPz6rwe32sd98GV/eYW7vSfSVJw/UEthqYO//NYZI/oE6KxPIUy/Z0LSAPTne
pviBNDvtsTC9bMPfzL8uRcq4EzjFUzjX8GqCvUzHwk3Tv0VQ4/2dfPx67WoG1opCEzawv7Pd4X76
3Wi6FPWzfYfvgBLOa0NNA1d8wQgWVYI9AqrXO1jwkmIHIuu4WE4p7+BZv4eYCFUdRrKHd44Po819
rCX+cKsc3aX11kPSyXcvQGgC9k02Xz2dBQHK23p3hne/uSvDt/l12d4bpTHjZ1oWQ1hgh1XZsuI4
tnRekVcFiAQQYOhilPLdn3aNJLuegFTja00hHvO322qKB7oIFsWVji7wyx6ndrqiCTRoXa8n7odI
jXFYhX9ZnpS6OTG/V0xxNwCyyQOIFXzsut93MJ2MkC4WrFPuzqui20GMOqBfmdfOGwLeRuLd/uPL
KEut2HTLksfATM3UW/iDrYj+iK0I+1TruXfMEG8ERVNFiPPcVWe0BMJ+AP36CxYONvE7wKJ6s9RU
r3GGi2zUVKv5X6tO4QGPrZc5j5uxuvvD88nubTi/EfSaCUA4aMDNE7BvUMhGIeGPj3OM6A2RPBOC
JxgYLfK4S07IwVKje/eyu+BmwAHAOvdOCVMWkGX0SAev3YW7ODKjjXy0qfN8KvJy6PEKIE9KaeMQ
Omz0uim19vuBMsAkCzYYJ+7eFHwwWKUDlE4HJvBIRuAp4QizqVvB4oIxN01bl38IDFjGKl+XE8Ng
sQ8bAV48rYsLwlhnfOjfErTYrvLFnMItQnH3+a9HIaKaDHw6Hus+WxXYZcuMgMBVponOChNxIvZe
HpB6g2O2fSka+C2PZhS7FyFG9AulxWE4yWn9oOQ46sl+SdA9VMPWKMKe2VJENSwHTgyi1yeegHK0
aIG2Na70cbVsbpojnoM7NnjHN+WIrLM61nnTS6kWNlAmnndu8VJ1ySEvHmbRn9r7nYLHH5HQrj5C
G22gcrAUpQ8mtl6sp4eOnq/lpGqvS42vqPNhO2PImqfxXDbt2g/9ElguJTdzH642jjqwLFB5Bou1
YNh6Lnr9kXQe9dru8P06yeMmh/TgvyNEoP9y68kFgi8O9Onmm1NyDKhfSlrNMEhf7Tv/rcOAFNnu
wxmFhoWpzTSUl+ZaJfwEnkcUxPC8p3ccbOKMfvIyfxWAx8MlmEBtFvn+FSN6p9hN7f70MUWpU6SM
ywPn1KHDpQNzvOXmQasL2gDvHcjgzu2C7apE7POEM3rTxlAVkIPXfj7C8BvZIb+22CJI3DlioIsB
LOHjsx7IWrkcHl/QIRSaY1/VTzXVibR4laaIcNXsKEOITPhy6Gk2aKbIriZ9McIKZvleywR35Wcc
RbIgWZaD/earfGX0EwEzbckOv1FE8sY5EyvLUftYsTZu8QHJ6jRbDZL+djca/Wi9sUJtZuW2gzwk
hGg7phTReQ2fGgAROR9LGMGtssJGH3HV8rvxHzsBKFSZar3Ub8S3D2dattdpwKWtxKezY34DGtiX
rPldxNREYax28sDiZa4dHvse9Kln0dF2ueouZJfXWNZQm2b3PzRV9cMsy1lCUv/Nf7DBEVKtSlWB
YVD449YhU6frB8fgxGlUPIAXUCjoggDNgHtfP5fmqW/mCXMMv8Q9DH1ie9PWK6N0UPGEbnjf1+by
xupdZ8yLx+CKgN+jB+Vl6ONls3P/31+PUzH3e/knXrtICC7vDOslZtOs6p1KN4cTxA6H10V0cIym
DD1UvsctFY114nbNgtnkR415y2O1WTx0C5KgLibkhpxa1z4ZvMd7eI9mRDef8wZ9KaQvw96Gc/6w
pOWE98bnkGhWWLLIroZv14Nb5phVQiiWGAAjyLQkPD/2/IrNYWhc4msCk9OJN9H3NdtwclzqmLdT
eXxAbWM5M/7ZKsCgJApYSn9gWDTxD6hE+AiYKTJAgjYA5aV/2OpCnk/MIJ63rxztpdqP35on0F9m
jP3wsZsIxmiEbTqaesogEBjafSe+aovBervMAnfaiv2KsDlQx4cFAWkHXXoksk+JsJh8rZJcNcuF
nM9+WLyYEgb7QHDUkEwmxOy3N1KZgBACvzyMbyOSrvOF4X9f4cZROSRT3cb/T/1f55g9TTj48UNE
MSjAjTmvLQESAP7Mivl01oAvBJV74CIHThtUQ+K3A6JP9KzxJ38+jxTjmbgKB6P0rYJoAq60VIea
KEkpLXJs/TiIQGxrv4wZvcXjdKjwMhWAqoDJH0CU6Pzjb6C+qq0PcdzrUv1lTCSLXCynU0APDESm
A8P1Zum/C55d2PE35HJQvH2uD1d1eUJRmLSjuetYUaw7K2wwnS5A8MOJvSXdiHyBYFY5ZRJgkbkN
EWy3bLMGV3p4SmruqjLVHxVGCjj5AU7nBWEB2c6YJ2DYwXRAsAnNMp7u024N5eT6QZumgrn7Sjv/
5sma0ufNbsBUNq/ZtULz+3sIKreEDwM5G3vAPlVIERM2ja4ccSgKzZhoqHjuPIm+NTffuM0bVMwV
uen/bK1RA160i0XQIUUYPQO3VJkARCWRVnd0qGxL5AH/81DtOQfC0Fh5Ea3ywXRS5G5780/jXggk
qw5gZI56E9zwqA7k3qdLS+biHrRABoj+Mvd/lFfADK+qfikqRaJ4qELjDS9KXdUdMNhp1+3rti2o
dv5SGz30JZamR3J3W9dRzO5uRtR0uVrAeldZDqFL1teBdxX3om8QjQfBgdGZTAUid3bhiNPeY3cR
Rdow67drmLvZstxVQQ068Y7NI8QSQXOcEY5EJ0qs9d5w9LEUQK4cxlMWLVsuZmAoJGoUbpJe09Dh
dKbni8/lgewNCPraQ+oniqeQnzvM73+p2FPtU/779TFtvbNtRP69qSXLiaqnl429GfadgN0UBiHP
B/O40UOhwO7slvj28B+tJ1OVpmnB9JVqX6dihUcPBqqR0H4CfLYiFa0RmqszVRVDfOPCY5WelJdE
cbD00ZFMIcNNWFQM6qDMP3esz6L5vqyuOWR27tfpBX4wbSjHSWcH+DT2GlA+i5CpIk3u7oo3/ibP
ozTKXDTlL/Rha/yRQ9OPUnqcTanscSeyR9RR2pYpMNkCbj3uT7EYgd4RO6gi26E9IR5CYaC9kols
j+3uoF1IXQpSsHOpohkytSx4UVYzwpv8XVUbKiloZr+d5vGj63NB5ItHnYnnzPf9AKgayii9KBIu
q95vdvW5U/8MKp5GyA93YSskV0qrRA9ASPWSBVnbw1u34P5foPOUie3uHgdzQ8XGd7Gg76cWZju3
6sPl7eKCqPp0euRpW00war2EwLaru9t14R88bb8Ssf7j3MegeX2Xi5QAzrmrURxBiPjC3rpsh06C
GJwZJZgao0Cm0hwckgzX8FHkcJhTiPWjzdOEU0/ltbEudDsW+kdd1cH0rIB+q396v9sugrRSYYZm
et/TV49te+Wz+lUB8jzc0ELeiCR355VjCEVxzVZVHxpYpb9UMtIUNpz+SL6L+vj0Qc3WPzjI417g
6hr/6Jo+zyrtRV+riYZf3UQ1TPZ71r66Us5ihzuMnPv58oquUzkNB40A5O24gC2rbNTOzpiNLc5M
DdEo7DinJODrS22gQNPSbRsU9MzMfSS7nmasAhFmYhCB7ybWt+xF+hVmY1LumPMYTZcSk6wDqVLB
4EF14BIIVSIjfyxLVUgwicbhUnqK9zvkggrrH9ohLJeFDJtXu89ARcLjhtd06M7b8rHmnWA2+hZr
aXcuvik5EBNxlpIGgfxjfhS/WyoLfz+kvANhGyNSdIdR/AJ4GPd8+Ky6a5sfD7FYXwoKMHqSv84K
QYp4MOXDaGMiF9A9st5ZJKslAKFYkRq3U2vPMgEtl5PLPRsXGoMydDyvfpj7tfe4QWgqmx2Whw/b
NcSjEChCew1pfkG1xJh70jJd3GO0lUd0nTkO38mritdj8vfVwXbyW/g2SfmqJMAZMTD6c9D9hDAi
u9zDv+aS9dUlGF3HJ8Sd7v9/ajnSeYKpAvmCV5XBjv/X9FhWkrN/sXOVI0J4kaMU9dXkFgaIC0nO
HPiOp1QjCE/EYUEawzomRtKqRGtqsS5FKY82yLLorH0PYEQiDv7SwGqiIubOKi2LYime6SB4ruwo
LKkCV2bxjahosGTwR+tL8CfZdga2lVyz/9BpXQNESjvblknI9gqa1QJl2Vn01Dx9achIX9x8uteP
RmFmJVnaJ8AQhgkull4Lvnj28y45tLBuIFvCXem5qaIEfXE1dmF7Nukwtl2WiaOcuvc5PO2zY1PL
2tPhtlasDPM16AsPNtJImKju164VocKZEqUnNs/aJqyklmwtaccdGnOOnoRIle/m7uQ8p4R6fa8Y
E56BVpjBVq9lrZrUljCkaHrD/W4NGRMQFczg+EShi+fh9qATgqoy1QqTcd0BpUE7W/VdVn1C6LH8
KsCgYDSxFiTm1s/aRxLRH0McLjKNsp4pwgMM6ssaZrvVXjbzurlNq1H/SBw3fD+F0DY31jOieUgU
q3I4WNIeQfUWnpMFQq3mD596RwV7FyPy+RVCIC9WaNdZp6d9jDp/9uJ8vShqo1Dr7L1NdFDKezsW
YtYiy9g823CAHI0o+amRGxBtmI570p6U7wwTVJijvnYN124ewQv9vO6tgHhjGmjZu+o0YQGQmCKW
ViXRZfvzVIVWW0smMzU7NZYIVDLY4HDomRZQGOJR1nFCIh1toRmUKzMv1R1gG7fg+oRWwdwnq23N
NUS0EKajNBVNNxJ2EfLOQYDkJdMIH7eKFsS49CS4Kw6C54cjQzmi4qq3CjB2bbEFEQp4TbTh/f6V
3imp7pwQOSkpk1nPmsM7rauKvcN0nlc2ikANyBY8QeYA1ZWwCbm1zhuljH+WEWO55XMdvp4gLwPL
r4A7wmVTyp21S4I2Pbw7jlUSEI30rZDrh3n9LaoU6mdjaCcctqJ+RYCk+3HqEGQSEN4kGt5jpLwy
UNXCQYFex+ytO2XfhR/TwMoGtbJouCmjO/WZv8Qktp0NR+XzbdJ6TEAM+D/x8D+0PwQ+T1mjZnqh
wmUGZgDHUC0unvf3PFZeas8ZjtikSW8iCB5hnBcCHMbpJN2vxN//1j7hvtTc0T2d8H4wr8qL/Uz+
GAm4t8qZY1ra24deYtW6SP/cpexQPb/z8G5jfrsknPYolO0gFv4/JeAq5RjIiMoe10h2jqrQSAM1
cijlO9UWrL2LaQhwUiadod/bWCrltcagsLYw2JBfCi9Gko/2Q3U3EcWFVqg8uaZ6zV2qRgSiscxP
QIQSEvqSfeGY1Ir193uIBNdD1P+F9T0MvOefc8DNPRiPsyCl0sAbQo75Ix2JrTZ+42lfY/vs5DDm
pFuX0o92jcXNrw8oLSA7tV6vyr6fNxQTLPC2/NBvF+mj7tNkuraURiNOgwe3ieOx3I7t8Rbi65vj
gB8C/SjZFiYGyKSf+yxv9J9Y89dxA7PPy/BYIbE6ZeIlEyFndNQdPKyctEm70W0KtPu8xGghX31v
owARlSUQz9PKL9ZP4DRV0uw2E26ff1HUplwFc8ikignh+z8iY1wqfLNdX9A2BnZrZ8CN71evaeZi
JPEtIkthsl+a+akZE4SO/ebakXEXAJpYW5Fv6iBxUwz6Qs+gnsL3yPQcPR4PhVQ5CxhtMMkowrXD
FrJTNQCvQVX3675xTIKRkHFmUeigb7Nbd6FlpcO/7RVjXL7tb54e86ydjeDQiHqY2MYXXkOSYZ49
GTTjzb+Ox+GZ+8FKWqF+/srj2c5bxHLyHbZPB88IUlqFNDJlIro9cNdbqXc0hO92FHORTq/jFdLK
uBPk0nzdAYyFnURQKTqgMDYRE6SgZD19p2rGJFZiuJVzxTabqWJPvR13JTteJkx+vZwFnwAHfOKg
lgfqiCqOBKO8mDQUbyVRUC6fBXlSbxXWHDlx8leGTr6dHtmCePbYPMjFzkCiRprfEHHdVQti46wF
wk+QSx4Pt1ZU9he8NqliNoKVo8aNaqib2fdvmA9yOhMrT4++C0Z36MTCjoIZdpf2njG1mjstaS1F
+Rt2HRLLQLmz8CW5GrYpb9JT0k2UrP+SADtD1K4mNZ4mviei7HTalhJEG29ougarA/bb4qK46I13
t31c2GKt3ur88xXCsKB6HaSzX1/Q/els6sgtCC3Z6qNNKnirnA1DjAXziLjyr+uIqJaRZU9CwQGx
lgFs57mKeCu2dqxryJ52QIvm+eOqjN3zhJOlGvHTJ6evE9K8xBgo2JxW7/9yURRhRYnYRS+Ouw/3
8BfjZ+dV70DAixk6eTf8jsq946Q1NxeB2rcoiH9sxfy/UxlzLv1NpCw8mveEzV7dnk1DizyCdPI5
0yop8nBdeozg4y3RT/Bm24rCCKnqJySaH1Pr+JaLOHF0FJDEN90KETz4sHxm6odYsNa6TXjhfeIJ
XBAM/IIkrn13pLs4wtrRzV+OeaFl1jPc2Fk7cSmZsq58qP5lUA79W9jBQdayJ6zFA8TPsZeJEWBS
DDZo/FZMTDigtjQcuj5WRe9Cn2u1hz/Z0x3N3V5NltMkY91O1oPMc0eH7tEfzH7LIjbNKflthDxo
OTvYzZXy8A7yp9Fvu5GagMvWaPOcSf/VmegSRL7ffZeJT7XM9lY9Rl3kxI7c5VruOlplcvwGMsLs
5KgEt8MAnh2Godpo2iAbo3Movq4pzHcdFUynN6PRFM48pMBfOjkOzObGgotI9fnd5hVKCdkcooL3
bKF11zYfXc2UgSP66xhaE6+ynh+jOwOe6/6jDZRIK8NNiFCHZ+oKeFZ4zQdu7C3mQRcEWk5oxHgb
eU34Crd7bbuZ5t7BA2uZEQINnd7UUGyg7MQSx+zLu2oliKdWIa+vFVh+UIdrJLh28qoaRcjqj4jy
6IRen8k2IfBrKM0LLxM80hbTVyVMfaH9IqKThuvf+6J8sQJA33ptOTIY/7G5ue0iDrrsuWwffkhI
5ZsJq3UPhQrvgvHoat1qZ2DWAtfujaZ4szhURocwGjX3gTZ+cg0Rv1merrYuJMMKOBOrZjgRyBIi
G4Ma1SNlH4w6AJoWEARMW1bGDZkv5Y+bPwoe9wU5gDka7CkkLXZ4Oj9IpkoIv5nSm4q79Q4OuMIr
DA0OaCVxqn3Xbxec3vbO5Rhsu4sjtLFQ3QvbRggk8rhKgieaoCmxwI1Yg0TmM4297kwHT5PSE1AB
JSkYSvJNu825Cay5d6pLI9ipWWyxsLKEwD3rjtMF7JZ7HHhnTyXoHP5AhUica12WKRnPtyKgJA+M
Og9Wn4rv39wzQ5WImOVB0TwwXMsjAqWqR+4Bxy9mCH2kz+hzerF4HeqI5H8YdmHxXfflEDz/B1Sh
z834NYqD21GomGEDYMimTsiGAObT6Po3npvsqLFx9cIAtaCWQxTnpG1a83aW6aI37aXnqebpF9UB
2yIbfyyOMD36BQCQ4r2SV0GICOIXC5GKt2y/hs68A6CaYAzEw9kYTK9irplD4S6kZ6uTHO9dr/UH
7IogbC3rRUAu2VIXWdHKU7escbTzgE1wqIifiY1893bxOhEJo7JqY3HsuA6HQFNhNKqRQJl11TFz
SEVtu0hmpzxK3Du5rVRAq26oI1R2sP/v97hTncVYr18gVVgi54ABt4ZFi/B72zTW/xcwp52vympM
5JPGj5dcrYavudKktIaqPUPMywm+uZeRWJfEmkgqBATFGpK0FkY/XT08Qje4wLauZIIGRz2vS9RB
TJQYNr9AdfVPFOsN8nKNeXO0Tiub0QXDNcoXCvcFSFbP2M4U9UKX8j8SraEl0xCYvdn6QRoq7spH
gSxZ8ECqhd7xkZXOuNZ6MJUb18jtTYwubQ6OOGykk1a47Im3k0XTTW5alyW+VppmhwYJ0gFtHW04
aOWo88UK+jQlpburINdx9ogfk+fD17wEtgMMJxBvMnIETduDUx80qdAQjEdLzmbxU7eg4yim2Mzb
3DwULhP9xkjaqOgCC/2GsU2QHk07fWoU1tGTuQSHVTWU/RM7KChccobX3sqJaHdaChyoyHIlnYvP
9ux4vLfN9UHvn8hfUbY7Bd01B7OHFoZojGLHrF4VQrP6hGkcnS03zvybEa3osj1QVZoXqghdDK2h
h6CEPjUwuxJgZZ2SRwM7ZD0m/pxMx4ZXMJd3tKidD7vomNhYwTIhGR2hNCb68vmuBTqRqLOaSWOo
16/Ninl3Vynxqt3xdV5msKIuWt/L1DrsX8XZJhbpxWbVzXSzQZvb3bTVJYkFv+ewDK6kQHMGbwv8
lBPobMyFIFAvanzjyN4rP5+l1OJRmZO10ewTXUfwXHToPV5JM8G7XvqDDzCrg3Dpb0uLQ7e1Or7X
sx/NpjzK5vkVHOy6O1sF9+3XaoD4PDxvk6PK7F8wWi7UDeiUx5z5pQKQJOyPwDJIMGgSSOo6Dltb
fI1mxQJxhJUC+F/zg8ic4DGc3vgdqzQSzNNca4a6LYdruV8lmSh2Rb5hDJT5rne2+PF1JN4ndNL8
jsouiFNZRoIKEhwEB5vVYBpw/dZzN17Hc2JZLRzF0XlKw9poKYcabmKq9+Qj0xraboZs4pl5sKnV
pVblRsICH5srIpU/HCzoi84aB5RErxnCoRzJnYFgE2BU+eUgVSLto7+uJzsmMGZZHeJysmllCy4y
WgOb1y6XzSshvhAmnOlz2Wy2W4UbLqfFt+V4UMsIVJaGBCJQVR3/S6Q6VFLp47aVxZB8aUvV7qCR
fu84TcPFx2v06eg3Y66kkUyattr8tB1gfRisT/VYlOmgfStRNq6t5K07pW+tKF0o6vuc0qRPvtiR
/B7jSB1XABZe6sLI0ZFd8EVQhyw6T1PgSa8pONMFoHCamwyb3BUbZsq9dhwolUm2DV7e7JxUE7r5
9Preh3ZJo+IEozyZ5dGQxxQa85q4pgQ8swRQIoxuhg4Cx5qUEBmhiMsHUvGY4CSZsF+L8AwkEfBz
9wKLUrRYjM8jQXxldRSLRROXUEneqD1FYJkt2eLRaTKuRzvA8anyEuxP3tE1zDHcY0RCp7bLeNwD
wV0Hij6VBH609Y8PGjHj95ukBNnDM2IGUsTwgRlDJcCO66QFqwtb2TPfhGReLaKhQQqUDUAjw3hK
320UfINBOsmChNZ6vrXcvRUkPurGJIZbSjsnHDDeuf/Jluft0KJdoPqRNf34t/KsKgh7nrC0S3Mg
ymYdeiKoXy7qR38JNW0QrDQNWjAz9rU0uWfltDo4VYWDNDwX8z9B6eXpeWTBzbkiAn4Pfc0WhQ59
dZZv5PGFO1n8+FmTraKroJMIP2rtidKhvVD78tZBCHC4FP6UhdTykEgb8CniE35pY5fEkY8ruiVe
tc1HXd0FYnEsdkqpVzfVTbp+dPF0zfGauve4km6Y0PsG+LXaltgqNjxx23Y6YFgCmk6kANfkNqvP
7vRn37FWlsQhxamYnaUJ4n3JxjHMtTHZ30V4uGNqj+fWt444iluDdqW9r1WT5C9RYip0hrO8SXRa
caY7FjtBiuXpn0lHqPAcEIY0Gj5m4KKKO8qOWgjYtDxmTuA5rcdWkTWyOGNgwZmbzL4eATFnVdhA
6kIZi9SAgl4QxhND0vKdDCOhviUhv/zaVE1fzUZYz6P7mWEZjm34xQ/qyjta8ZMqR9urvZvThmd9
crDZpkVribYWMD888AzT4/8P107Dz8kUYXu9jA5dXJBLqwxIhTgipcm5tq3I7aIqeg+OOBi6kt/b
DdettIi8zwWNZe9fQ98Y/45vFFQlci/ELu0pJaFVuW/SsuyhtdpyiwD/p3T/DhamjciNy/zuu9ig
g/+56tLKh4Z/4KzCD7CkUOPn6ybHGvmfWGjV8YxdFxTLoDjSmae6KyypLBeeb3wFHheGduLMdh+a
GVH+h3pDISjhseOs2aHkvNfLKxyB4QJpNBTwD5kHdXuVZE3aApmYlARoqc1k+8Kv+e0wC2VF2ef9
yEfpxaectkmQEuSApIsMpgL110W8c5aLdZNAHT8rowKAP3DO6QHRtrWJB0X0QKoWohEogpfNM5xE
mzN+stia2SIp03lTFw2+Nl8oTeFPv4tQ7C9H8az+TRbV2wJKwWHkbmHQQDA/pYLw9zYW6BKfz7zR
IEoyYQUsy4DyUmRMR+QTfuWnxzpmV4f56Q5zMV0gY36lmb0zItujBW7bRVS3F4tNRHmQh3ke+/5S
ScnyAQX7PTWlbtdaxudpC3IIESkhh2yV3rpKVjbtVfCxVrjgptPXDSeok9U9JmCzWfCcqHo7p0VY
vbaCEi5b7nEE/ypiBKHdNdxrIZePwuQDre1ofkGO2H3HFKkd14Mu328Q+Mh1cAiLHabuWPiBy+uZ
v29dQVrhmDhmItPJMgMwBTz2uE+IdSkRlTtvHL+6Im8wpPRJI6d7Dr1+SSyZA5EGPq6TwMMWAIw2
6d71RcKm+kf+2hAu20VIsxRICDyXh+NJ4Dlhto5Ry2INCJipHVwWFGyTjia/FVV/pPm566UTuSIe
YHjOseyyG6Iqg/88ywhLVdeGYj+iok5VtxlabSbaBvchLNAdLgJK3DE07CCLJ0EwiSyoTFf+ZchT
GexBzb8IYoGFlfjDIrp4cifKdyisTwhT5UAjjRb4WmHuWBWGYlXa8TxwtxXAG3KqH5LVrVjKwhDr
EC5Z9FCquqzJ6AP4+sSIsXDqo+X3ND62p9HGcd3G0R3cnS+qULf8RTL4NOgwS0tJ8FU03kUVpjmd
EJzclUAVz8bVsWiiyx2NpFi+XvFd+CrNQ68tSCXzjAjiIhn73911a/SHtpKUmJs3+5DrvdNah/aU
OHnoRN7ExCRzO9+aHKL0YiNkUrZnk0jfN3AHvsbUDTtcow2A3yO/WtV11hXSi0aicueiKdExbp5j
4GxjsydKOzX57j1H6kBfp8jVdqh6q26Ao10GCmJnb8MqMhYGifa+LGXXuW+aBTLTP87wz/P9Bw2Y
VXpqGRdZug+uWbPkMoHZUOo8utUPwM+1t83sb3eP3bccMREnYotA0cYrv8pUQN2vuMTk0H9qMcpQ
Vf23utN1K6bS/bnlgf9UQRB3Fblci+0IYbljxNdqaSnnFKHpPgMJqhQzIp5jDJ0bVkXOprpD0NaP
1TvgCzHPBAPOFqHaP+iuYZz+iaY4e1qtY7LLws4Ki7630gepHtE43tCZQ270T74rOBRMRsXy+F3J
8S59iGX99umB/Zt50adWnKD/zwIFs2T6MVTN9HOveU0vURBJzgqQKIChlBMeheGtsL1HDFELOkqF
34bpKm1y71MpRgGYqUgHz4G5maBzpXCBWynUJkpuQy8EYds7rGidYfY9CDxcgF9SMiuXqLrTy82j
RrFSqJcX392+6JF2NcKKSC8HwB5wZGwtDeoTpVBdIjgAwqsF1RIW1MAEDj+XMm3zEW10Zp1SWInS
n3CyeZ0VfFL7fYtA22cuYfbPFSrmcdFJRLRddY7/Lnrg7ENySFPUaFIEsI838VlhSDiIe9PTuIPO
yClAiCBTduMgU+F3Y1LqY3GHY4NrqWheuWk8HPmPppTumqjMZTGV8Xj6HoVMUvw7iM4kaVKQIrj2
8hcRzGH3AG8IW7PlnRuc1Vuk7TarMWOUJ/R9pvp8D56emG+4RuOMozpH53KPGFoXh3CKp1Hcsbbx
lGOXENfGhRAOeBaZYKx7RTA+hrWA/XzceyPYLtDbPAel7i9V82/EvPi2Qm02zRoaTwyLZkEhKFfr
FsebmyXfaS1oOcVOx8E2iurIqXGTuZTMx/YDfwbSX9U1C3gSK8J6hDZWk0t70EjvY41MPyoaH/PL
7jcTC98FoeeVpdob+qp0L2GHsZF4X9AXxXYH/i6HUQmIKB/jmSAUmwCx2MeHlznSiQhMujI47bNq
/HFaIb4CokzJ6UT48N6rXpNe2DY915v4TSkyjIYpAEw8v6Bs5QDrnKUVp015b4OkN614hT+ysCyU
VQjah05xkoI5yRN20WVYn23PWrhzEc57XXEFSlz+RDQsnb8F4LQFjzBJFTiAD48py7Vu3nuy9Vfd
bstea3U735aBbEkCvHKJ9GADbdPq2onaU9g11QMl4k0iL+VFduKBRlb7PRHlPBaUkPVgm7F1xCAr
+RkFpDNnpipbaxyLGB+VD1/H9QNnHmLqIdRjGOvPDv09wIr3lM1DWx8cBuxtgEnM7WBTonvf983f
y87mCCTcb9OZ7LR1fru587gWWi4iUgTFdmMjhB2zNuM89LAuaFjHB8a7MbOX+QxDc7/+9HQAFuXG
e0KxiTxJvFjvXVfxniQq2STyOVY1CChnYs4NTxsJmt2iQUAJRIbwcA07jVehFCObRj4riX+EKWZx
HfX5Y06F5I/8U+zSXZA2AWqtke4QvussZRhG9R9ukViRVr+J6+iWpFW7dS8GoklKruhUWGJOWInP
FtAqAg5749rAUs+qPtrxyWqnmAwBAYoWSKzU2Q+It+eUT0+jCTLz2EOsEoYtznWWlSBNmw2Q5STG
7a+5Bp0KnZL51T+qldhTgwI4B80+Wue/N52W0/hVN/NwpzP3DnYjsq9yDFf4lFTMvinVSn/DSyxx
KQ44mXj8nJ/AAe0KrmFnVcp/iMfoPWgoLp268KwDwpXd89Fb3ziYrYWPSGkDRCvacSHn8eqeDdL9
M6QBIueyasGV4riJ69uEBvFrCIN+eAn/KQT301U4MvOQA+fhKbc60pooIhvjWEf62ucZuZDSUhxO
3ww7gWjFK4Uw9TmvSQ9F4k0exZK1jCa3yyKmWKGnbZniSNj3m/2J9quNynutYtUV70DN5uSgmHby
a3Wi8yroK8H8OUF6W7fyXIjZSUfTl4bTYlxPvPP9gtE/nFoyigdvIvg1CINVVUCCe8zMlSPJD4Hj
egKj9K4M1ghLsNInX9mM+Zw74JEomiln971TBmidkNdfGHm56e35Yq3k/Hpt8rTP3MqUoX6KOYSc
JBXdqDIiLRnSLxKA3GST7m7pCfAsDqxnh/otNrW9iPPZ2dBcClEYKIbLeLbBvcxd3BTlxNvnehCb
pIsnsL+1gluBrycE/kyDPlY3Hb6nCeUFDgtp9A1qYnql7JFIsEEc7ZjoprPvmaHg+yC52fo5WkDE
QY4QPbB60bFww6MkFQzRa0kKd3nVtTQ/fmpsWfY7SCCTC7PbaN7D8sXyMtJ61szJuD9Pa7v0FIFJ
NllxPO+uN5nORc9Y/4VEdounQxPQx+w9fINhAF9yCJIjplOKxTL42GVAcBQ+wioeq5F2I44jRB/E
dgPc2K3wRfB96t37LPM0jOGF6cyv8YGUJGYVDlU4yJGmDwv4EpWuciJkpacZ8aU+p6XEzPxjCuOX
R5F1vwiytrUklC32Rm+dMLeqHso36WgRLKbIUdd/KH0bIM53vrqxAATSSvaLE046NgDD2dFd2i3X
nxPtwbdiWQKweYwFP7buHAOXqJGW/XiKQI2LAVmeqbuoXKDUlYz9tXWAzbB2VFXEOwMeq4UWM7s4
VylNszXBoPaSUMoWRTP7DfPqWnE8CmVUZr9+Ld8q5x7wbJcJxyzsNIoqHW9EF5PzjesXgV2HFoYs
fCcUpRVnosrwo8ShfOB+HoNj2JNWQ3BJt1LxXcq/XFjujmkV0KF2iqwaOgZTmazaVWqAPC6JAcAh
IbnfDKvgLlb1JkcQUqSCghmCxpecAFLvn6bjVPHJgWsVZjX0k6zymL9/seC0oZeLHRsQYXXhaTVY
O5NZtjZVoj+aTji+7IeJ0TT//5ydWZtEw+t4fIpe3NVDLCnlOgVcCdXxcmFsHUlUZ3moY0jKc2+b
xbQstTrPPMCYSrF5nNrn8eK9z+7goLFAOOz3Hlwd4Jct4iOmXQr5+FeomTWCaXMbNUjwkSiCaK/j
3Rf7XPoaQA1PB5cr/eaPB/m70QORmnxhh3974OSWsbcxbRqvh3QYQmHq2KJtxycZMoHl1/tMDDgx
sAJjMxXrXHxJfG2rDgoGE3ocSKZ45TMffzhBLp6URcQVHQZni6mvmRFK8KpLKkqwBT5fu+PTSNqt
xdGs/B2tnmK5t2Rr3oVGIus+bB51ur7hU4mXa2onhpSbuMFf+CTWoF8y0J1HqEqA0jA5HnKLk3VW
feaL/dggmWlYsK+jMpy7PFpm/A2LIJ67X/smKrIJ/1lKvOa2e7eRpUhH7LmR3W+3MA6G43q1heeD
t1lD2oPOSyNwlNQUX6CMuJ1Lg2s5GoBVA3p8IbJDnyQZERzj/EP60ZgwXiwGd7aYz3EIpi7vurTi
INrdZyJpBBzQxSL0eU2jHzqrkEqQ7710+BQqrZrKZakcJsb7phXaxZQ9H/82rMn8yAdeKl1qAXFk
+IOFG4OVa1pw9CvHb3M5/IgID3oJIa5+lJXcJKAsSF1uh61tU7zBW0K/HtxM7Xp+WiZ3m32wluMY
fbsdctDhQ5opYdqtGkghJ8SnsITMMc33YhIH30/lVheX0WPA0XHhc2dZHeq9GdydUibC4JfuE6n4
zcY3JxLXqdwj5YCIJAAfuQ6ab6DDkihOkxyEl6QT+bXo0n1S2FrzFQi6R7ewNiAMMVGpE09QrAw8
9UJnS4u0L8o6gPX4+OG+daZzLAwD1fybgj+4QNwK6c3DvJi7RxM1NYKiFkyntHfRd+i65/xTtDjY
uAK7KdxFrWZk8FTS+rFQMBz7YXWlJ/HbIvZo+4i+LHJ8gChbABAj0vTv3j3x1pxnvlNmDzOrH4BN
e0HMHtPCb7bJ9faV/APYCTwuVqZFnuI2x7dahEaZCMZH9xNfmrkC83nRdycwHTZ815ufxPWsh0bu
nMMq3AJvThcLzmZsaRyGPFhAiadiHO1yLgJmhPy9K6UoB21rUmrXgaJ4Sc7A5xAaWjemdYaMMNup
W8ksLJ3OXgK/1DLx0H54HWIfuJW7xMFJNjv+vCnKy6iHqe1PENhNtegTEcNsTQD+Dz0EwdtZIMqq
sw52nUBmw7W4nsEGsITkg5WNd7N39GGJ1gNlHfSZr6vdAUwRe18VPXr4XdvbiMYPDvplbTsGUbsS
5JC0TaS0q2XS9Szvk0vDvYzDY62QPmy+pL3qGGVsh6ViF1m02ZHe77Z+h/vk8k5L8MG3FL85jHTq
XSPnTd0X2cJTMO19g2z2xyNBVF7JuShxtk7Q9ZF+m4oaCEgfCLGanENXBp3PUeqQGp1jty7GSnSr
shYkmx/pYDQEGhOavVyjr2R65cUDmJnD8EMQsjA7ctZiSTnZz/nEyDnvUUoH3MDvu8G1iK+wurVW
3Gg2Pm4qXxt7Tu+7cXoojHm2ggmJ4JOvpZj5UqBrk7wmm4qW5dVAG7UBY06mYJf45uMsrnKgQjXW
Y2HzXZL+VNu80wvAt+qjwjLOwXV6uQEGoaCm35ndt3gdgNnq9EJr1KvV74gLaPT9u1rYR+7TlZ8E
vBVKOjZ3Jc4OThPpM9lz3vVce1pO5s5AEDniuChZSjljYXkkLvunytbzU0Hq5FRsVU3ZWPgSfNo7
gAeBhV2uhZ8fnML5hQyHLGoSe2WSKsAKMmT2iIpGhFG6FspysHG8wWvvh4icRiPJcHUXWyscsN3q
WEBxqWFiR9qwUAK0GAkU1V2E/rZTwW8bSItdwTJmgNMQa4kPVcczpp7NjU/IHS9y92ju/H3m0pKB
qpQC2VpLvPNqC5brz0qa0KVEmvPzjk80BXhZ3rptMRUujkPWadzyL0St4NDHWIR44p0btQGgQhgp
aIV0hw8GJXfB0NUFnm6gGreMppb+N5gdadRV+27eqVVx6P+dmJx9KTRqnOBw6s0AgaLuy7tNYoE/
4ssqc4k1BcZIJlEXf0RxAOJ8O0GepWpPs8ONzbDj1h2UuluNTtXFlRqalebFzaevt4fKvUVDwVSp
u6krAJUlx9M/ttsW/ZTPFuID5Y6vq5XMEf5ZpfDjh9GQvHS1aGOTHT3CmEwCmv668NJyCV+vzHBA
nW2XP/01VvRqJHjPj825KKKBXeEPeWsoqhFUpGwF1rN+pnzn1TuXCf/HCL8agxMUc5KNfi7yctXS
mRtyI6efLmfWJo9e1Ego4xSVd6GCDDnR2JLf4AcB8YAXiYiWcMIQDgXa5evLQ0F7MeYpY9xCiK68
1wUZlH6KJJqFyOIFAOHm+UZKZqGljdJZ92UpkOfau8MW/ghOWOdcPu6TouLnhVHnmX5SqT5Qedfr
KaS/xve9ZEXFgzFRzHXTXMRNx2qPGwGRAB872CtN8Ibe0i42g7Y7PJ/0KBZ8ztUIVdU7/d6Swrnq
ZwgtpYZWY8gmiXVycrJaiQ6v+vPDHuI7vJ5nDtMGo5TJRVEARPPYotsilSHdxIhEimA1z2Ed7Nz2
CjhMIMXGF/i+lDIioD3fKO9gdHgea4Op9gNlYmIvDLjavmshD27m9TlqerdmY72i/OojUXwIY9OZ
rz+d85Sq0hjACXMyefthaM0uy5Zo5YDRJwfCq63E8XcMg/jx+P4HtNGJ1z4xi5PlgzLWqSFEgt77
OocEfQJLGS1/k7ctyifIhSZvRo7ND1q+JOcEmErioNKV+/ZSEyMZsQwuMwVQVPdNtXCJpT2eHHQj
fORrYcV63XiEJq2+wUXcYVP9sxcUNoQ6giZOzKvQvDPq3noEie1FMFokFvM4gs9T8Gv1ynp7PmyD
CAPzoKxB4n0BX19CLWRmpG24NluVOt+v73xjWqKP2FOs9CkHYE/nb+8RvI2C7Ww9P23HAiUgjoSl
1warfdZ5/laXoVL5xGwp/HYV/awPhGeFJdnctxdwdun3k1jpZmZnWyaE4NxSVRbziHSh2DrhKXxM
Pk91OP0Gf12QufUG5fIUtwgh0J7UAq07ua8eZzqwIu0GnlV5K+jtVD2OYYLyjdHCl2R9whtnQ4nF
ICuOr2ejpRRPP46rbxa3c6peJ2fF+kQ05oGawdXGtu9ueE6hHXyP2dP2++2Yy+SmUe0OFyWTm3Kp
QB7KV5I3h2cfaRG6SsCk6zXdBhOVpr7A/hIlDOkRSDg3HiJKX1lLI/2DTFNfYCRo9AfGEjoj/YVI
blGnWSwy0P402fSHiWpccKdg7Dfzu8ODYyDUELKD++N5cliMmymPQbYODQrvoSoLobY/al4/gS0+
yW2gcOH0Ke/VLeoING1l/YVxv/gAIhCQ526RsUOJwo+6FQAHuhjTlHDee1pBZuQyVX9xYNqlhCzO
0n7q2nuSY2629dukzMteA2/aHFFoMpa2wV0GUs3S1vsPI5ClU6Ys18ojoLN/eRR0LVv9Zf85krOl
b+jkCHSf29jB4HEMZCTRJQOkimzNvhUF1JBzVeHw6B75jqYiMKfTlXNaZNOoVsiYcsfBxhtSOjFT
qeNHVa2RgxgSKbpfzqxPcKTsQii4sT74AsnMWAHCrcCF8zzQi3oUxmpNE3iGyqjrfmJ6CzxynFiU
S4OUy23lus5LnVzq9f/8DRmvpS5oLvEm4NfU/qs0N5y5dpzt8zmtLNZGiROjI6LIfGE0NIqkKKpr
BPVrqbkdfTglq/bMaebZ5Nckv5KDAZ5Cp1HBxUCWB2VUSECdkURgB1SpllHZrMHm3pNDt5HgcDoT
GxlGoLsh/dX827RzBOjwGUzIuOjr3EKryKuEy8YA3nF9f23xW+xKxuK27VjngPsToX01/pnaYvrE
20hlSv76WXC05zy6TWv80Ss9YKkcNClgwb5FDBawo2kjE9mwVBDLnamEMcKx/VrayiUuHiOiNpfz
Z9mKT2xKGyk6pCfhi4Q2RrD2oicqaeJ/qe3eMPT5+RmL2esz68rdQp2YgIsvz5beu5tdu8OiAF0m
XnLj7Syy3rsn35ZwcgsGjun/zpt/hzCnYoW+hu0pARXJrPRUc4kAqL7zURWxTqQkJgbUoDH+lF9Y
t5e+ZZDLQdSnee+baD7m89YQRgZRVSJzHnbTmbGN6ffhQM7tA3GMArJfssMXTBCPtFTCYEOaFoZE
vgzRhhmbFFXuFQvg8SEQIjRBxyzSZqpFxfNx5+/rF5Pwc4Zt1iuN6nsgzmS9Taq+d7RNDIYXP1Jr
5VSo9CH3oyWm8srDPolHrnMN2zaSFL4RRc+hekD4yOtFmU+Trg8vSprRkWtpeQLc8Vm0ATgJHmwu
ytWq8Pd4PV5q//n+Z0Rqn0BcALK7c8VG1XUzyOlmOO2Of0HOeehXjn3+K2LPj/BaDtxt2GETAAWd
I4T9Qa3cA7LQbdmw7vDaOqzt7AC2XuTmCZtzCGFNf4gCn7aOuyRJVu3SAhHoAo10CXkNLHQR3Jaf
w9Hu95jqdn1jcoYZKrIrCMsrZj42GcBumdpF9ZgMidCb6MGwsowiOZ23XDC8/XIKzg8fCpC4wgKV
wiHlwfswOTjNK+8ky0s4DClXd9Ooc6Om63JMm1DLjc+Mmh6mwV/XYZ5OX4Q9NgYM1iVvynXJEpXk
YuFpIGoXQiUY9arSl66nOEQ4yfqUupkVX6RwBgTUsdL7t8fBz6Sn7vUhc/Gt54XE7q7vB5UQizeL
Q9o3598EBSJeJPFVtenIa8TRPpaqYRV2f1rKlmskVZXJNUPuTOAKA6on1Bo1G/4e635++pgz901c
DA7DJcq94+1Y5fzZ9TYVwNzGjniMgo2tG4c152nzBsDQmQmRFQ3LJmkKJ4EYKhZ0Ou9xCfhCreJ+
0bGrnJF4OdC/9/nz9kciZlt7ykA2HG1A6jOVOiwypFzUdL0Htd3PIitEOXbEEic+2ToDa2+KGgTE
hglSODgJiQfDuKPXw63NCzF7qgJrRuU2Mnt3JlyJxEu7cLIwbCU2cKTB76lfnfFAdDZWb+KiMOD2
xJBUu770I8uAhcLSAPnmXL91q0+IK07nugqUpbQl9z3uyG7uHzJ43iOgmuOypoyB2r0OGEuCgg8O
+byG0KtFG9q15YUc2994EBlQIN/z9JHoZA98uMMonscdbRJJ8M5yy9E96U8YQrLJGIlkCjRB6gPz
0eR3CHR0pfFAf7gd5NTlvNXPazvlZ+7YzyFy68uu4m9pcbira5pzdkhOq2gwDk1ewu71lEEs4RfB
b/uxu87YVgcjw84ywRMjC7/I3mZC8imA1bwyyC7aSFbLsLKrjW26UwF0mGMgBVSn0K2FFjf/UT++
Nd2DgJ4VbYGafZ3MzJBSkdR0XDH+3wtcy0SQNrooAtY3tnriF+S/WUX1UlMGuwx5kgdhK/f3U9rK
sVh57YtVtorIy+Rt9y1i/DpManPzUdJ6XzNMqSbGYqDZmtToooCrt7W/VNbPmUikXgIVEaEaiNd/
eOHLmaC/VZqh/RC3+sPaKg74m7hgoUIScwGdDsrf1rzcnC5UYPpFLYZgzKPao9rpOFQLcwlOI046
VmVCXk96dwS64V2WD5ubKO7jYp3KCjY6catVJ1JeSQuXqEMPRbkrLdxlyXJtrGNP7tF61f73ZyAg
AGNuKqnlBThgzhIlTrtBxus5rpsiSTjPLoxO0/RvzFQ+KHyQQVEMo7z4TTsYPe7pcLjEIJ3jwx5U
KIMgnnrqdJmH6MDbyuSuMd/OlQ+DHKASac2fn468t4lxMZmXBS4MzIWUTlCeEReiEDt+97aU66vy
32lSbmhbEL180M6YnLL47nAqLJYj3MskUKaIUhMmz3URbqHeKCAGM1VfrSfbEPIj7YBWgSd5WUyU
ijdkDQIEYY/hDrHqiv2d/KJ3/EidOqKjQ4eq6F1TGrHEMIyxiALojHPrKTLM0PeVmiNiJ9o4k5Hc
8rIQK3307Gw/UxRHmJ4igo+wYMbxKBJGxTxDocVySE3fgjWOJxWpoh2gnUJD0lVlFEmuqE2jFrm9
B5rTCZ2hr5rnJJf/Xmeaa1dkGhuUh7dYzOd6qyAq+3CR2bG4Zquoo0RYqBx2jM34bxhShHcvdZQF
ownTqFLMYJVugYPNfa55RLFeL/Vk6VXBX3FdaJJ10Lq6PSPWEfMMnorx99cMOA5U/5VFQlda99PI
PpAnKLRpCjqF7wshS5H6V1kTKym8bfPdHCgR2olZg7xONlhrFGkKCBM2HGJShAo7k0rgfAzfTBz5
KYZZE2Dmccvd8lkOQ7qvtcbXJYpGNc2sdrEqNWO2o0ofdryp/KjbYL3FzARm+zzrlsV1GioRhLwm
fmdQrl1kEnhH8dI5yq8pz1plqUDG70HfncwNIROxnJm+bqMK748wyYsE0+pQpr1X+3RUq1bU4uuX
vaqFK36rHahNUuaWVjI897YYWsaYRDSdeQgGr3kVqO8PC2JLN5vFVIe7OzwHa+y2OVFL4L7Ql5IV
Xj4VcLW2E/4gzdpvl/NKR4vXbQ59QThX95gcYdJp2LY6w0O9Q+kBrKYIM2ThYp4Kd9mTPWnEHDN4
iU/VbvovxayE385ZZGQbuNGE/NzG249ztu6gbJcuCaNiIBJJPoHINgBgAwvywRmiNg8iWh/eU5Zk
KLAMVLJiJJsjw26S/EJFAOg3CZ0Xiq+PSa7RxqH1a2rQwCGXLj3cONptkeq1yx7hN47s/W+2Kzb2
+hDM3aEJLv19xabw9bl87DcHFPvJZpqVpDy5LmO1tzPKjIdWjY+y2MRxGwwKa5hkT2vLBS93ARZR
XE5Q7Z3AFRcM9x+IPwMR2jfaMhcbiMWl0b5rHllJWsrcYeBUkxiahOcs4VNu87UUh1zioXAs5uar
NY5WqQbiCp6hDUtRhaE7pGlZsMhCbNAoiKiFp+NxkHlkVJ3vOgFUgpHa0Ayc3OlkngffCa1vKtwc
cKAopI4oAl1jVCmaCu6fBcqWnKi672FxCDy+66/OImj58phGZGZ4Edg1vL0FQqbWWE4HL5Jlm2hY
b01LVJCoFFJG5h8zaR5VA7vornGViwlbNeWEWRjAoLg3So8GZGBUth8xbzr7ocB2amsRGUPcs0JV
QnXkZ8wNtRLkh8PnwudfuSFSiwoaob/R8kYz75q31CNzp22XsgNdVSckvXEXAvjX2ycm/hL8psbg
8xPtzlv696EtgwwqFmnsGJBotURbZXI3P/RoZn1Q8gmJAOBQ2zFKCIB5T3qhtGhPWghUgDMMOIj2
9e/O/pwVF95T+xW08GVBOcpC3yBSMnUin6+c3YlixLU20aE0vgu/EmxViaYwyDA0Kx0sgC7A+bIc
QTtA0hPsGie20PgRedU5NomZOnMyGJuKZKdS5TlQDMvEZHEDfmRweeoqzZzIPyN/KdlaS/dhwBFG
3bFiAOZHzKNA82PiHpx3bU2r2u+HSKRUiLJ1cnAV8d27LxJqHfFv0RlBMef4RqZXGSGgP9MVKt+n
blhdUAvxTRYjj2N67b+9GE+iaTG5yYEs1HHr8T9R1IjWeKGFINHx85HSZWOcO7J37INYBzEDgBlN
/gMc87lGGyLuP3j40WvJhiSYH7HJCCPAYL2st3dVQVrVr4PDgjGhDnudymPiqsWvmzQlYUP+CuzD
jnP2sN1cFm1oIXsVi9a5wBv+ql5d+S8PcU3hLcvNUg2AnInrQVrG4G0FG7GaJPjmXMpP7gYoH9I6
ynLnK1ZjPjnPrsSBzCfAA/RB4pABVDJBkekWkMZPYQ/wScvrsCml4CVqH7q4ahvv9VS/9e4wNANW
vrXW7Zi7zXs+Cjf9YG0FVS4KY1GJA353zZJp1QT/U2PR9oKyreldgci2k7dna8IV4GuIRyQkJx+B
FHQ0aVMB/aAy8xok5iv0SWUJ4Rc4k/jyI+zvGwqu2zEK8MzVl8klMP7M9bhMKFKR4WIKBwgd+xSk
OviXDMhQJ4/NliRNWq9Hg+LSZ26CEYIHdN43hKGtRbOUaGLFOdxzk4fnLK0YKPsomETF57E22rco
7lmDeHx5FeBfYX9zoSdO0wzjdHtioZ+jcAS/7Wx3cjpjlE4K4axUbk/h5bVTta+LOBPXmjCCQGBy
VgFeD8LmmOsqKm4eQYCl2VXBMvwSbdOjZnLf5OfaElx6GdktIGLXwyjdsxSXmUlFH5u3cb5gVpS+
Nrh18LW5VZlUQVYotNglNVZksp99Mo2IeOoHRmOXirGaIOekrixpRX7dlnfnBqxtQBjiBKIcMDGv
cuMl3T6gc44vGoPCCZqxX9/ul+8/s+1hd9pTP0NXdcK74vfnmqBqQZ15PIZDCm4Y9xQ5DOs3NhF1
wcjn2QwceSROc3nvt0oTTL38l1wVMvT6tPiMMces2YR5AEpp+G2hAhhO4jOQgP+DKLI7H6Wv+1mJ
mYmzUqt4T7On4TbQlbogUQsg0SV4GCfQzzyyO3lIcuq6THs0u8WH3l8c51sj0INKFFUILjxIdHwh
ahLHvKY2ZP9r6Ne/lPNOWdj7v6FJd0KN+nfYKLeO3b0tRDN/xfgDK4UQ+v0HUKPsaioNKwfiQuen
qsaR0O6QBmjHmCIdSaR0fK/sO8KJdcc9v6aAn/dmRLFf+KVfvujFby0NyzhN6IZjUj+HQxn0/sT5
rsd3WjpPKhhY7Ab5JHi4BLo5p0FjvMXoIXv3C62qT4KplKeGG8qbxAZzHdt9EDfx/PFRWEXTQfwl
sCUpXb+k6soemoZJj2RCKJsxuPIv9gbKXgVl23CKaa4sfBpE2x6fgLpu2igLln+9FFYyPZJilD4s
5XC9ayytcUrjfyYXcdhO9IpN6bOthOHbXbe0jIEBHG94N2q8nGn7wsjGY5+CQuTO5Eq64J731riZ
mmB0ZZZvimFwm6GXAabSD/+peyferN4462hbiyXk3NvghUt2RcbOQ9GoxONyGStl5KXza3Suozkf
O8HKkAww0/TptsOvGeo/WX2ppZ5kPrbTr3eCuSAbKZFbTPtqth9Ym8ZkF7CLiCa/KamIC1e2YlYF
fV2V2ha6RiD3+W7t7JagH+21f7lc/am0QwGUrWmXWCsTf24iHFCmNYEmoppNL3l8ofeY/npruPcP
+X0wKCoeFm/0I2x0Xnd8LjNcgbZ5sxy4pCIVrMPT5Uc/0yvk/FlTSjj5mbtdScRi/sKZUfjRE0rH
Q/vjcg8ot2/oxvSwcedKEcKRM5vLxdOxPwa5irRqlLHxx87JvvZ7NB/wlBZEkZ5WCm5EWm9bY4Z+
/PLLKQgT0nhy7ZyVHGfN9KXzxHY/ifIalFyly8FJVxfEnOGzTixUNU1Sh8RR0V40g0HO9TmBhNaR
47mGQ3IltOlg7j8abNGr53qw7Dejm7R58lqubJ22A9E++craKFwWgdTy/wzYYvbCYvrP6o42cVYn
Pba0elknf1EF0+Ao8IdrUqvgtoz+Eg/ATQtg6tW8jOx4W0qwQS3XkNS0m6bsSvEvLjvISx0TVDJP
l7liiKVxfdOLgeaXpXDsYyfSIpy3PtJrJIkM9I0tLEEPS2DCv+krRfVxET5+TLcPysLd+XuEMsXo
TTSRUHOSZmwuYzxg9vyObKkPqro43sCobSeiVDLzluyC6En3RUPPDu5djBzRy4Gm/PZ1ahKiWUXE
I0ZScD0EAHmfGxkSlbDqfw+nWWMO6Eh0/IrYPaxe2457iWQCvecXkb0V7mk12tNooZfT4orplNlo
ywh/FHA3lLIvMwG4UMQVspmzlJRI9rYQMAm57ZOU4Kv7djgklC4NueZ4B5bdf8JgI0Qrwr905pj/
MZN9GAQEVftoV8jOZVZWcaeyjiKSod1iCdKTb5g1MEuArpBN/B3Oxmg3s+h36k0wTKVRZYLaaptq
Ov/Q9Izk/rPMwkZfVaQuXyqYH/8OM47nfOmCmfmM4HO/X8YNdFvUb5tjntB2fUyKybp90j5YPjWf
fKEDFNinXa1S1JcMEYga4KdlACkiLAIQoPoASyKZEClHw50A/ivmF/Mkc8CVP7vXt2GBoNADXV48
D04Mlvl8ywItfl/jR8OUtiV9Y1aSTicMq66IWFGrEEQsZVefE/DqxlQYCnII1EVtK/gItrBqQ3uC
Bjbv3mJ/zPi9tMnRgCD48zzpOUuHU23pCu1Lh+obmBDxOJdmV6SHDpua85FHslHT1AcM4/+EmtZi
/XFS4UzM8/EAif3I/c3HAxQ32Sz3ukAVkrOzEx57oYpGb/H0WVYFmrmhzBN+zUFfOU/zLiHLJeNI
+CRPCCouoFw+WwqTDrX0wS2A0t152ok01sMGCJwX3YjUFsptXaL258DIRrXYZvFRzgTleuge/S/s
XB1r1XTYueUXhCSaEX0f04xyDJLHjTaP4Ix9nkKNJPFLdX4aWJHCZLu12gqG4H3vXX0Isazgrkfb
FXiWPE5XcnO6T7T/6EnvSXz74c/87thDXD+DovvqoyWbmp5FM7o9VlixZ9PVnPe6OGRVM+oGor1D
fIJ2/fDm4XOQv25iGy1CeNZXhSAnWKl7saJOjgTs/qTWfJx43BdpJeQaavlCdfD53FhgjyKnGp/I
jjaJXf2j2CPoPcgtdv8c1+nxkQMwqSROeNRXr0C/mmy1Hj0vq4+BqUrl6BNy/MKBTVRJNlnh7rGx
Tnsp0UhACy0cS0m02q0IWgcrFdM2zHoYPQwHeFzojs6Ppf/1dzHcYGcKDPgw1t0ZsEJtXKpMr63s
3Dn1hefP83KAqaJtYd4/uWSHvsNgjGeujNTPHQaONU3CG7qxpObJMSR3oRf4M4TJ6bFAfERIPEno
vjjqydon8UyYEsJ3cThndPeNWUoalB0G0cxfNIz5udHNrDtqLWfrFvn2lt3JUAqKq9sBpndZJAfh
5iShIu2TGxPClJhUwwykXZq5XbQE927k782sCSSOvV9C9X2bLUil5EWNcm3yyYVFVFq+LgV3rODs
3f/AuhMPUjqYJD2QVIy0wL6/D9AmbpVq5REIn1pl9e9GSp+jtteie/TyqYG+ZTWBj8JvfZjVnZDF
W1f4tDK7iRNTWNBNZJympbBU2PlxNErnguEpbrm/9aCkBCpEjdYhWm63NBoFTUKH1NfgJU9uJuQQ
oFlKAl+S11Wd2jp2WUOc62T7ywFUuhQnQOiTR65AF1V/qLd2PrGL7bAy6ZRzzimaVG+Vr3iWNcv7
I7iiK6KLvQhcGbGI2XhabEOKSvKUMHyYzic/Uae7fQ5EiA9GFEDazNdoO8ucXV5viMgXveivLqs8
SmKKLAS0tGegoAJMY88vz3c9GKsTz5vEuvavbe8Hf+MqNUNjKvvUa5VsaeI2bDKoIh0f0OrDABiO
UmdK6UpW9h29Jus5B74tDFPXD4kanEcrKelOxSuvo061j28y8OQVNo6zM12hRYCVpyBzyT+hDzF+
En+J5Iud+9L0TKFY00tMl+5Shx4aGBiN47ATW0qDkubjC4g5YHrNpmfhEeJxjlKsFb+nW7zWz+wZ
XdjKentGeeWXYb6MNVbwRLxgRTRPJZKe5mQRQaz0sElLXmG2ZkxbEwt1bS1uvXAmJyrg8itqttAE
GrYrdea1FXggxyaooRYazYF33KwHooL5OK4ZEsJvc5/rvFC3/wlN3ioN7uDz+XLgT2hgi3USA627
ec3dfthWV9Z1c/eDn3OTIZ73InJ7WEa6H1OJasLqFqrq+RLaCC7MAnVwKWDVbp8mNmwlF8cP0shW
9R8bXVUF595UjgK2KpZ2aWSVLHQt4mGvkMZ9qX1PpvT+W1qkW5fvJKnDn3U9J4BMKGccRZc76N9K
61zxyOan7dGFtgBCO+a0syfzRqu+iagRsf8MoJLn9g4+wLXNmus6XA7jeQ1LajKCyyoL37n4HwBz
VP/1SXfZgAXGs0/wTBB3ECmVdTcP6Zt9ZWwJ5uPK2zu3I9WfbPnFIT7LIeGP8X9W3otZf9AZS0Wb
RQBpPAzOoLiWAMop3djE1GXRYD9FaCqgK+jlAQrSpXL8HMOW3ZOh/tIc674MUn5LknVRWdvBWLUI
99XaN2f5P37Zf7sAitGEBVeA8Vgb3C+NJkcfTiwDHogCXK8LSOpWv7lC4pAMP9f1ZzDDItnoiwWF
aEw7lPHTcj1KLOk0whGDsDBPk3b7TgmVcYR/fzCmoZ4Zuq7XkoLVmKcDgf/yK3cK0G92m1QqE1gx
hGFEu5fufIlqTh9p7lelNt95wkkAT8iXf4efX79O6aehyPDWOzJspMmxkpPYKxqRek9I2+qfTP5Q
VagpJ2qJ0KpkM7awafx1De6hph8DCIpmXVac2IqiYqm6a7/moH7wz35VVfSP0eZdGY5cMBuX9mI0
t35D1xApnacm2kNAYAhA4xwL+ABnBbalcUY6VFXwq1w87AO9kz4ajPQrmVXIIBDEWshH7bbKWngT
ewgOJ1Mbk1Wv/3cswUIiljzJWCzCCc5UH0OpdXBy34SIInC8KLpQqI2idvSqvIn26f3JEV/8DyYl
vkkoup1RbEJPwW7gK0Cn3PGZa0gNDF3/zPp0tEvh0h7jt2s54Cz3fKBMGdsrP0j4TIOgjQvCRG10
GbaV06XTFjFc70OxRoqu16KTyFq3oitE60dLA46o39vFkUr/ZiucITcMWdvw5vf8skOV1zpVZ+S2
p2e1K71FD/1tKi7TMmQdNzfINpNq/Hzh+cYJ3LS81cJc3SLiqEek7MhYjR+6ZPHTRW8ENAdnn64b
R9AzdokCHPaCYnXw2Z1P3lfziOeribRtjm9q7kxlGh8WPg6xwukDdhX3zr4gLHRuakWd1K8Pas3X
KcgaHKvuXB551mObLfiX5ZDZTIkPT/Nqaoi0h1erdm2HW7I6VeoixGwhOAnPmoZDx7xHeDHC5skb
sfKt1lcBHcAsdZ03kfz5pO0n9IqIhr5D0JMAyURfoMMiPNeLDYZ042j8FbvPi32Mzr7KHrxp5p0X
iUQa163S0HjrcrkcrhHjAvfssrl1bBu/ah+I7/hwo0RYxEXn67FSA4onkFCo/4b47ZMZpxmhou1p
Yvf1+8M7CcEitA8wJw9z2iBZFH4wihIuX+o06jYCMqAVXvH1gBpQF3GPaOQ0uZvQDDE7tROxQ31w
n98c1N6KxUpR0CnmcL1FPMom0TE6kg7SDFyfA4aQppdagZN5HXId6QAPq25IbXDDDpnSYItL8CEB
lrbusRVLT7ZoUHyDxrQyr+tB4Z7wycHa9rl+Cr3RHGh00gSEtAibjE+J8lb+IJ/plSfh9uTTnEu1
rFpsGHyL8QSpZuny1g/2JHzzDtelbint84mAe6MRO/jx2VDYLQ3KNgZSrbpw2H/6cdiJYjSft76h
2RqvXcn2J51ypkO5tHH6FRYu3kyCFWGSyA7z5Al9L7frbCQbv0pksWo3InqIxzO4PF2VeIgksHn1
tPubbrgRZijLGms5G/0pCZlLCv3zkJMtzY0buachx7Stku0rmApgEc26vc6WXFN/mCg//IY8eWJN
Md8mriCZJSDOk4bvU+eXHl54bHJNk/6WOcYxIhsx1ZF5cgnG/+NaAnb2GdJOQ6jSAEnt15ZZrSE2
SpbWA7Jbtbb7pCJBm9l11WS+Gfw63/tv6deA9bAiLslzE5DehgEm9K52GUibHDSWS1KccesQnb3h
s6k4AZmi6CrEKuPAPLOAgBS6MYUG+iSeWgo69I8VPo609+PHZrgQkIoasssvrIyPmodvLz2F/8IE
RlV8UyOSIzDElNS4nh0LitF2K8aDz9wqQCbMc0s4Yj2qwpiZ1EfY3yaEtMWAVeJRynndAVsfR5Pq
3X333XQOlpBfP19W4Sz3s9MQBlmP1tS/I9lxtJjWkEpB2wJXp6tyvT+pc8IyXkkkKJgTdJCWgJl6
0NzWGunNDhzg6wlOtuxFN1b69BMEpIh5r2SiHrqv/FI5ttt1+bkzmJTyXjk7+6FMZgVpgTF/IhjG
YQ/lQ5+Cv+20S0D7Z0TswSRhUC3qrOrni1QemoDhFGE3SyhGof6/bIXXVE7nCp50x/1PCiADtTST
edt1VYH3HkBzvSvWL5YYW990Sgup5c1YMrZC3iWqpneYzEQhU+xYHsGhoPigehziU6ZVSvgt8vdI
2ESQVw1R6RRmzBFRLwroOzkJm8J9jL46DFe5wytmc6r82jvroir6yFg4re9u779HHI6we0SKqRTM
a2/bR+FR7frEu3Zi33CbBGSowdeOmtHikVp8Q0DV/7GsoH9VylB/2qISv5FDI4gvg+FfEolkja6A
1loG2HUKWjSyv3iAZEPz3GN7JHKHj0b6eJZ/ISiqHqUgTQC2xdlYu9SDuWHKt3WZTauL1J9SUgys
1VzxqtlM30OO1qaZMWaG04/TpMDwCQs/7BtLn3p1TpAZl/Gcsxx2uQJmKZpgPIL8F26kPpvqVgp5
ynKIZ/z1haLpvLLm0FW4dmLpj1vg/EsOtqjdRovgnNitkdf5+00rW+vqjiVuTbFlmOOYZwErydpW
FmYpHWpAw9SxwCmQkwTqVYoqkC5iijC9UnnoLVhmpP/MYVK7tEkaLKfxr+Spf5/GT9gEb7vyHvPU
O1nLMa9xHvMdBj9ui4xqNIQYvMDZmuog7rHnMU2qwcVLb2OnxlRqUVOSP8nyYzHOytJ2Nfz9vQ/+
IvZjYA10tB1zLUwub9REZoNjvRC+2f3dSc31f5BOfs2GIGSmeyNBXbzS633IfiGHfv9+srRSwR4Z
DyP0xKQtg/mA78+c8yOJnx/NLQB3kOYc8iWXt2z9OWn2ZK75klxmkKsqemWKJ/em314Fp8U0TvrP
GZhvJdA1tfD5+9O9aZbXTD9nS7QkZP86Ly2zZKDp69UfnkiYRD1UKprOYRHyT2tTEJcjkM+iJL/d
zoiFa0EDMu6PjYm/hKlndaJQ6jZ4ruPp5rCAsY+WoGW8OFpDluEJLEt84bKZ4P+fuVevC8iQCdXt
s4/7MhvchclYDz2OmMuFTs6baaUc2rkktNZ7iLgKJaRFgJKa/hrYYD2Zt2K9ZDqqeYSFcm9aGoHs
UTKSufp8UhWo9EdoNMSe3KKjkxY58BaoY8i5g6FSipVxRyaJN6E9iek+oaPKZld1NomhePCEk/Pl
D/2FeF6jjszpYq7PuhOS1OPRAOnCqzKU4I9ICosnH1JGUbqOGO1U/kdrMiAH09AOnOazoVoadQNx
dHs+EMW1i6bG4Qdr8Z8FjbIPVoQtaA9uPiSvKlcZYNbAkcjPL80Ymlv1ntRnOexsFZ5HffW85ig5
QPKSe8xbybdpWP1vZT7kr0WIU6I3UoCPuGnXf0znx+nn5vj9f5tkoHfNGips06FJ8dU//cGzR36I
LZfVKp2bnvn/fNuKQ6348UJb6J7j9ToHyJfPenVzQjnY1GMf+qtDwpQ4BXqembD43l1MKOAV6N6b
M5WPMOWYl9Wax9yB8BHSuUe/mbIaN6oV78iC9wwoNvVRKKovUySXUR83JdMSelG1stGwyyuvOVRu
GFSPi7W5HwqTsJbJjlMtvbci1021621NwdkO1w1J6Ig2w6yhS6XqFHs+cmsAqbOMuBww1XwBWX4J
jvQe
`protect end_protected
