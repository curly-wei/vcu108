`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hH+7Of7V0HrZN7akhr/PGWzFYMFZ/Rw1Y0MdJHcXbDfy25bCrbSAgiAHzjAOItzVH0GJHC0TwaAh
l8lQ6Djj5A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AmHoZR7VmEL3tVmWsOV6IVQew/VOu2KAm4f6KJfAzXGRTTxsXlPXI5eOmXy0OQc+dTQXlc4Nyebk
WOd+g7avEM/H0dDmrnyrAy4xkmGgWvy/yoSRg2NcrorlzU30DXGyLUL7cC0fGGT3+aYDfpalxOxG
vMlnYmB3ol3sAa02k/0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quTe40cgTFzwGZ4hh0czXTRPjRM65yQ2xuoMk4KWhGRBXqG0mDC0qybq0KDkzMvHMO9o13XXh86J
3lmXd5z2U8qbCCQTiQ5D5fs/vDyxOt2D8yzeP9Nz3v9pLob1z25U2A3IDkfdMys+0lSQ2Kic2K7X
M9l4gP8XjJ7XaZMV90LT+K3emy6GtwfHL1RmLLmz0wvq+4goCsSl98hEr1onaBQ9FjjXJSgHTEoZ
asLa6XQpuzHvUdrr7uow2fs6n/v6lPMa2QIEVAOBRHRZfcfQ8mCrRActebecw4kgaKOLxGzIWyFi
VJjLlE6Keg/yDxLLEGAzIe0fXmz5IeT0hi9g5Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e0IXUCRiGRcDhitPNE5pcnOQjcFm6XyOGSyf5ehAs8DfcUjdAyC39hcyh7lelM2n1wk5DOyQUYdV
sH1HD1x890dqy0Bm+/WUTKfxQ5I0MfCdzTLMWpdnX0TYkOpM7Yw8f7rYC6qJM3409nB55jo5jbXs
BAEUxqIp85fdzNw1bsDtj4/QyVBwF3hP7nFhpQv+EKdvqv8Q0w3KT9MgfmK+tlzpA7nQq1DUqyYL
tY84oCcSfcuA/mVkkAZzSZD+v/Q3sdnagb4fc0bpcJT5TQnRzdluhqgGQtVo9Hv3B/rAkJ133atf
AhgpSKBM/HuMkZ/NgBMJ7PD7eVL6yIU2qjgBTw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h5kgqPrm/ghas5o50sQF7CkRrd0UW9+3Bgyf9II/ObYHKU5WTqvdQVx37RiV6Zuwx7jY8BKGUrC1
6GljDBL3LJhoaR694OorSigRqGQq9DlbWwvPpubN73/pUcAA/BmXyPJ11iAur9DDz8dL8u0AIVBZ
JMEcSp98XKgEOnXtjaU55MTSv0JNClbz/1GbpUB/la5GmUUPVd9VERL915SygcAxXa4efzVDfNQe
TDR9Cg+V+hNwUsZ4AL0NwCpeNAD+IBeM7wr73ySKSUjSInxlA30lGKpFr4nZ6c/01uzl+nrIAdot
iHHtG6uFhJXK84C4UUrX6PN4AXNBi1ScXRAvVg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qMPgyiJBLpyBHm6njnuRl+5NmZjHACVWOf0ME8HZlaAMEUuZ00geWO2DJ0BCcg6vVw2jNUSHe2YL
wAuBLQt46RfOun3ifJd0vZ0OhmxMdGpmaBkF+pDreoI/Y+6zbpN9NLfWQkPSbXW405FftA6mC0LY
RxeVKPNt7taRM3Dn7tk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GOYJBmvSniPrLCFEvUHh6c8XRUg3Opfv+CEOXcm6o+imohXua80ifxh90luGWez6hJmfSTaDELfP
EFF5QnNkriODMphgc0hRiy06hmsvCugkY/+lnM1+vmLXcLsYksCkRp1yvno838j5TK13b7OUrqjF
fpYN4rWrOt+Od0qedbEyjVw1DaVbqvMeSEy09YrquzpAB1Gn42zQnRqbZyB3P7UxKxd6Je78SneY
ZTMyCwaU8UpZ4qBnHHuRlhiw5mnZoM9BogaBHysLvo7BZaDOif/Zebq6qPrmHuj0Z7B8J4XLLpKP
kYrrZxtmMkKcHsR8kM8j5XlIL2/TVXXoecYL8g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QmPcEzlUpwA8HkI5E7k3BJ8/+g51Sr0bTjftiABHZ12feKb0yyUwc3DGo4XhaK2hwP9A/eEaRoma
DGsRKeLWw0e3ct2vRi8ep6WFdF7j/Iem/cY4NZlDwWOsU5p/5aUY6JIjthh9yRXtopvvMjCYzfsJ
/aV9biiKpCoceP7BX9BA/fsNJMkN6Uz53KSeUPzAHhAjmqbPrq1tftbyHQAdeTBIITSgKrbeoJwD
MluQlsoQv6FFc/AG8Xo3Jw0Xz2SIjACi5gXO0Om2I4nU923OlhwwBiwNqVm2ItyIp8VbqOkoT31n
b3utr1501a+m4vRbYf1P+coW4adHWojl7PGtnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 4944)
`protect data_block
iDYfqNwlpRopY+1YWynzvdDiz4ihvWKObGnB/CbpM0ndy3b8HYKHOYVxW73eYKS8P37UZXFbZaRn
OswUg1hlZrPhTv+I3noV7716GA6XzOsL1/Hbb8a/r+QSTiBjM1cmMUbpNDNCiFH2M932r/Y09xqc
/V73QHn3A7mj+1vGZc2/J4BNd3fdF4t1vmVFS4VW+JMfRy6bdlmZbGDsJeP8aeDeSld1x5VHDIpm
TzaVxzIoZAlVpOEaWFsV2icqpxNFgpXaqIUpARVBRYeQAIfw+QoLWJR7ZZ2HNkWVxrGqbh6o6Ib7
vmdAAithMBK6yPa5sVj8yPkao4DSqVGslgdRlTGu3HgYnVRe6vdJHDuklWQFpFfqo+y8ahWdVIEB
x9qxlS6FgB9/54xN5wP+mx+BF4/DENE+TSiZDYDd4FulfUKPv0f9gOrs7r2WD3XPMNwVl/bETqRP
ZDPs90HgH/jZZOaUWOv9HzyDs8/mshvj+nvuw4WZjG3tQWjwu7Df4XOv8nrdyCU255NP6LtxtCkC
sDeqhm1paAM69WHAB4++pgHSE0lKDOmJ9HxgPW8ik1Zs58BZR9tAAmYAjbDpgC/yNEDcNGoAzVcY
k187W5flT8N72DfKA0rHUaFhK9vCv0VPdiEZYPFyo2a0Bmo060//1TzXHmdRjVwcvB/UoR+e4kzN
qjIdR+KIlqcxJMVKLxVcEL3At7os60oeOzpDv00DRvHpboM5L9gMNVG+IT7sWLwNnwJvNODS0lLp
8UbL1jDOHzvcn/WkizcHvszO/tu56RgDUT1Diu+65b+YXy3D4X6G305USyEGKOLHP11cXADvMhHs
UuFwY+kXRrL021g/8oatOmWcJcErBm9BcshI+ScLlgbx0+JmwGhQij4OFJi3svThoxYYxcCr7jKR
PqBF8hcMvxAtvd+oIY87ooiIaV9Wl7A3yOwOsGR5jK+bpdg/lwZb6nK4n47PvEhUSyexi2DqHFRK
IeYNiKa8uB9gmFCmWqcBbjn69JEJX3QbFxj7OHbR0piFY7ZQA0fY5B7cmrO3xbXzUGUPlU6J2gBS
Dg2J/vMsYr/CyyD5/f7D2u+tntNMm6an3zezaOlm065EFGwS8I5KYPnlG1xStHjNYsizIGFhPD9Q
atGUEA4uxIr3/qE9xqW0qubfNmwZYM0VHz0kzHQt/TF8XvuHg6F1U1MYZjvC1r7Z1C0MYQeThLUi
NXB612hprcknVQCoLtAGxTiBLePR2wBcJWUIZD4EcdV+OTx2Qw7Nz4zbGXU3RePeEMHftLxSmeED
HAdbc+9ik/DQG57uEjwX7Rvt1JZLS+QEUlcnokOJt9W/xmBy3imwuLn6PuuhDjXnz99ZK/JR/LLc
zdISxjMmnF7SvOpjc8k7DIwvCPilnwYZZFBCXbOw7sSzg+qMCUNY2kpU/Es02eDj50p/7kXuKpb2
qIxPK5qY2iVUe7MyghDwgAhfdudbei5uYycTaV074F5XWlKU01wsOL6OqNYQoC2OtC01Ur5nCOSq
Kqez69yRYnr7WtSjn3GoawfZJuy8XNtoNoP0xIRMvVaQxOO62Qcd2hDQKdjr2TZIz6+qN4n+oN/4
Do9iQT6C7yjuaY5kfHvXNgBONDVM1b6unOvtRi7A47fye5WAZNsJKlaNf7x8b0Hkn60Jsvct76g/
IVJlSpL1aExl1YokKH1MnbkY2vank3ibJefmfv3OrkesVafhJGSJfsrWKUWcgZf1h2kbizwuE0jz
tEuwnHIXfD5vmabMqb0UgRFZh7TCgPCscoZl96Z74Y7cnIamq3KCamMb4qBsZluUdZOVVLhkZ8+W
z6ARwODUBLpMg/hzWDPQSAb1NEM7ZSFOMtsbkE3DmptQgxrzsOUvaA1G77tKIHXkeyajlsovRNG1
Wyq7aZpx7++7tqmRQjVAGiiqiuNAav5tr1AxrqSORwHjN7s30vPG7/VQfKmlwH2m6NSmrxUiHHPF
VcxRztPn+o0PVpiBbWDLQkzjnA8bi79yh5ESnKQWJFv7GP0hs834ta/Y58YazHrNuBuzlr0nuID6
FZI7iXUjkqwS1+7VNDSwhWqklG3wT9YySHSWZc3dWCM/PQkSskqH8fjpgwMF3Bphhley43Np3oUn
Hzt/xrzYemmUNOR4hUK+L15X/aKYRo2fyJ5UjcK3stgg7UCFgYuqXOmMxjleVvLIe4C1q7B4wh4O
AtbI1HJWPGFdetN+ZguMbWjnI04ALdWch3h6lZQGfDN5jiCx12fPWoFNJgt4xXNeqgcrtsyCLvIC
AlCim/SXRQv+UqiQ7jwbp8xZB4xcL+ELHn88nlcskFNbZ2AN73+AFTIdmanDt3oa2PlE6Tpu9fkz
5NEElOfFvxtFsUhX21bsCeWMYORD26DEAdto91DQhLYY7t5z+vpVudjVQsKUFpXyi1iGCd7paKAK
PA3pECnxEpDVfjApLyCGoRRKemhnrPFmvclCl0Q2tkuys97boYFHrwQVn4LFXMrT08RDktJ5Ce5n
L6bU2ZSqCk8EWSOYpxIXP6h/zJpp6Kh0MolfuKlr9oMxENGTcW7H+dmd+OOxZn+nWhKfV1uzSXMu
UEiIaTVc/sT8L4fm5VT4m33h54cG/kAXjTZrFQo+iZnOgkXRSZF9V+X+o6KpQCXNrVkSGWCUTdBu
c71vzwIoswEVUOrvc0a+zZvo0qulkcghpNBdG6EYNt9PGLzim6fvhzKPNE0pigPvQQMPp9kTzsdx
MJYClbzqedj6ggrtyG6XNDzfAYXwayAeSuPelw3HH10WgyCthQoKji3WlfzlB5Wq2Yv7J77Xse1b
BKkBF6P4jCDxbEcu07OG0xdmGAEMxQ0gLTQYW7+Gf9ybEDH3xYEWfife5XU83ulKxa+reoa9w78e
DL577szLqi/TkKxjeCTG/6YaN7/pqPRwH2operqWTB087NIfUi0lvKrolr12RPTaf3aehWaUv1Px
kdlNGawkkM40KyoIT89c/8kZop/fJFyJcM/yoGjjvnTVvhoYsrJQxHFABR6BEB8JzTMDu+jV1ByN
xysOD+O2Q0qJUxMfj7MLFPXAERc6/nW7t/8foYTNsLsdOcMnrn31qHitT6VrYf0tCtKgVoIBRmbU
ln6GBKZHSOJj5IgcNQ0u4keZ+NBHlE3PCbV2QK7H7FPhRhwC9JmBqOzIoFMg9UZYfDoiA4irWD+b
0jqjfa16gQ60YMuGc3ApYlZRs8TxYtXKFjGwQVLUKIspiO6jpIRyuMSkuy9Mnuz4cWTmFVXmKPDu
8p/ytAZsRttEmATa4HqNs18TUqdawbBR3Sbw0kc+Ow+H4S46XHYyA6WTsBEbXiZMvmQUn56zdjAS
S4MTZC3I17og7p0Kt0ObWC3NkQ7jT8baLDL7deioNXMkVuVl2P/UwR+1PHN80Z4K+eFfrXBgM78r
zlHiRTlvVoxEtbnZMrPaO7J9prNZEWzSGKWuotkX0ACimF8qUYk4nb6O6kEdEhmVmSQxqjiYbi/9
5te//5jQERJsUcCv4B5Ez9EQL73ajyDk49Gcy8PXpzzht7yNglaWwJOIvhOT5ZIi0LRjOvoJXaim
+2KDG7TGl/pc9Q1Zd67sVw/U3Vmd7dyG6FOkAR5zSMKMfBnKi5DBNHYKQqB2hOWX7JKc7yuttccY
rbw8UpNQzeOs1cfU/0Tg3FQVzMzMKH9hDXJ+YBjwovXP7FuTL0vQ3Mvv+qWp16GYL4rTjsieJi0f
XFAxSiLFA9NBqrAuupdHCimAAch11atHiNWr25LLg9k9uZPshStqMBCPUuAyQUa/yAoj7dWyC2GV
4rICx0aDioQX7WEWmTt2bqtnlMRwyHIPPvUFnYA4jX30FkGZLlYmwBVMBuk80np8fGx8S/Oz84EA
/V4k2zRNIljk3J3n8k/w839sJaEnN9wEL+BSo28frs98rStI4aOHMqqXfAG7qzFk/eIDkMgv0WXa
9l9liJYfzsqOAnqJ3bQ/ZN8m915fvqh2mUJlodXJ3FLrbo50lLXXoplWCJkLy55SHwySGbwqNfXg
TD+HDOXqIR527ru2RytnM2wgvVZ3Sxh3vzsFBa9iizs884cilKN4/u2UOjfK1DeJGEgTGZvyqBnW
G07yoshLMpjt8ideiCrtGzCckNxWcXqxrVQpZ0s7hMJzXUeetEkgs9qArDfzRAskylXqd5LoGiaj
42cImo/o/FlJrkhd2Nni+R/UkCkr2TILQTO/OE4E8vw18EPzGYx+7Jy43iabj3HJ70WM6KHDX6sw
T2BlWNYZ2ne6pU9gFw0If4jR+jVVo9QPfvBspP8awq3PbNfAq58RxO3Q1hJFwnuUzkqpY4ZLT3If
pRRpUW+cNTg780ABK+5Y9hMQwZHAwlgdcMU+0dEcxz75Nk1fEM0z276zzXmCi5qnCbZOepSYop3M
/Ulwwr4ryWCpqxcBDHKqdMVp+J8qlUBoDOR/cdfxEDwXbVIXVFYKigrq0y5+B/ItzRdgQbaje7vZ
emGiaUSkfajEmO2veSDUbfHes+PonftaURvXfAUU4puM0D8f2TrYfywWpjf9qAKzkMOS6pTq6ucR
8BfeQX9ZprUt93GFNdQffqDGlzGVwLwPah7yzht3tfkCJXbMbEDxnInrZUetjQt0eG1n+NiNk2e7
G2QtIM5Ye4VZIEVeAX/90ItUsw0SUdhsqTj8741x8Oq2i8PSRqbOxv9n9PmCpnO0Wm4hNXI0mP+2
mhGkj8SPGNH9eccBZQT+iamqtCvKhG38Ku9WG7x3DIaiMOGu3svJW+gDyaRh8qAM03OcQslzVm+M
xI2p1In3kl/V3U7X34pQvBGZY7gu0bJDfj/I50PZadyCsGdQsBXj09Cj3tRFKI6G1eChRRO+ebDs
5ZdDg/eMKSA5tQfKiHNAQlc18wHtiOQcRrusTHj5LbFD+F5nE/eGpmiM9NkbFS1qXyps77me7ybM
Vr2SNmaqX6i74IHqJGQYdDEcg5GQ7HxkJBkI229wLJqBIgQxpzSYHl+n2TwGwmjRhni6MGQw1qP8
kIVW3WQ3uZEGaa8sOLYKWYDTW8uYa1sT4k1zLCkgzOK0N6R3xvsfgpdwWcO8WpgSUnqMWEXp1wzs
CFW/b/Sz3XByYb4XxQffbNt0VSert4Bf7x672s3Mz7jpl9VgzfErVd4ShXHkfHLAjXl0WXF++oLT
xsA8ao4iSF7xb+bd7bdtNO+SNSJSmNeBKIH/6up4yHUF12Fm8VmRdrsGZhlhY/pWggquAUiPIYxF
KlnXzVOAmUOMIEgiryDk5SdRpaxNaZK9QnE5mZiwksvqvNed6Fxf3HeQv2y8J6HVsSjRasEj+In8
9ASQ7TaBrrZAIMB3BxoZHzlcF4FShgRvERaB4AwifF8BMDxfUKPr3WyM0prFG8k9egQA/1oF24J3
iu9/KC2TkqD59G3q8nTUVzxU0kF2Dxky1FZ+olaxHI7S2gCMMOdfVGjiRBk02MyLBCWmoNkJnP+3
KeFIYOhO5v2rmYqEwbx+pDlEIOvS/dEcf+PAAhO4Cm5Cxi8w+F01w+KqXld2G7UZe+MNtkFh36Tf
EWT9lBoZ5l/uxKOhFcNBmGM0N09vgSLVR8XLUiSCt13hBhxCUfoZZQg2rMBRBgmwOECr6pFVucan
K9x4nm9rufgXIsUuJFxzM7USeDXSaeNQM36GEojwZAFbQrKS+z7yBk5hEFGAETG0z0qd0CdtMjVt
5BgjXHrd2gv/Ku1JuDrTD9/rk4TIfUg0p97SKHVU86Q0KangZyvNY99aBOMrmwVqkHXdaNFBRcOL
uhOY7bA6hVFbtW1nfEgsq+244uq5otnZgGRsBq2s7lVqQNonhL7KsCDI7QdpYBGaNdaxb51/usqq
TVBY96CraPrjt3XEya6xwjcSBU6e0bZTYV0mxSvfrsj+ISkESH9Se9gdG5rFi8gi7lM9SK0UjS4Y
NTyQdN+1xaMxzUjFvJS4/RUmyvvUcZsKX14phENuWqJL180BP1BKTjglrIDk/VKQR3Oj87xjiVKM
LHu0vB3eUbNaJRNGtupt5KRTMcuVlLHvbBydaNs0WOhUUQLEEzx2BhzpTqVLWhZP7n1lENta1VUp
RmcCMWWEsUrhxDCAL9lJXILgRuqJPhdvFxHblIn1MCHJKJxjJNh85bL6yiQgSO3vZQIkt5JoRdM5
kpeelWVLznpRQKqvFDBj5+p3Ny9EdW3p6MPXvBcGT5ROqYl9sC64OcwNHI9hZxU033lCjKSwuiZD
Owp/SDcfyGwSRSe2mBknAA0K26tpCFQJfdqF+yPKbwIqFMA5d+9L9u4LIEQp19XDYpi06FnWMRnw
u3y86LzRBU1HpEJc4WDFFEwlf0kXx4npkt6W+Z3v+5/o/6QqjCmhQgW74EAqKNkbNAs72HOnGt/b
zwwXmz5i/k5VtEbcjNWYzNYnwjXq7xW2QdhVbLVoGdaDbsqrtKMA4ft0zX82a7d5XLpYrTLBwArP
dWurfEgf3T1t+FPtuKJVAq+8pJkPe2q86v9iRPa5QOI71ozoTr8OLX4bYjy0gPaKu0CfPHGQVTCV
IOFMTdLSxUgA63z8IYhF2a7sys4gVUcv0reRM9UtanUNDKth761xdKY2
`protect end_protected
