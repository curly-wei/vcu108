`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hH+7Of7V0HrZN7akhr/PGWzFYMFZ/Rw1Y0MdJHcXbDfy25bCrbSAgiAHzjAOItzVH0GJHC0TwaAh
l8lQ6Djj5A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AmHoZR7VmEL3tVmWsOV6IVQew/VOu2KAm4f6KJfAzXGRTTxsXlPXI5eOmXy0OQc+dTQXlc4Nyebk
WOd+g7avEM/H0dDmrnyrAy4xkmGgWvy/yoSRg2NcrorlzU30DXGyLUL7cC0fGGT3+aYDfpalxOxG
vMlnYmB3ol3sAa02k/0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quTe40cgTFzwGZ4hh0czXTRPjRM65yQ2xuoMk4KWhGRBXqG0mDC0qybq0KDkzMvHMO9o13XXh86J
3lmXd5z2U8qbCCQTiQ5D5fs/vDyxOt2D8yzeP9Nz3v9pLob1z25U2A3IDkfdMys+0lSQ2Kic2K7X
M9l4gP8XjJ7XaZMV90LT+K3emy6GtwfHL1RmLLmz0wvq+4goCsSl98hEr1onaBQ9FjjXJSgHTEoZ
asLa6XQpuzHvUdrr7uow2fs6n/v6lPMa2QIEVAOBRHRZfcfQ8mCrRActebecw4kgaKOLxGzIWyFi
VJjLlE6Keg/yDxLLEGAzIe0fXmz5IeT0hi9g5Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e0IXUCRiGRcDhitPNE5pcnOQjcFm6XyOGSyf5ehAs8DfcUjdAyC39hcyh7lelM2n1wk5DOyQUYdV
sH1HD1x890dqy0Bm+/WUTKfxQ5I0MfCdzTLMWpdnX0TYkOpM7Yw8f7rYC6qJM3409nB55jo5jbXs
BAEUxqIp85fdzNw1bsDtj4/QyVBwF3hP7nFhpQv+EKdvqv8Q0w3KT9MgfmK+tlzpA7nQq1DUqyYL
tY84oCcSfcuA/mVkkAZzSZD+v/Q3sdnagb4fc0bpcJT5TQnRzdluhqgGQtVo9Hv3B/rAkJ133atf
AhgpSKBM/HuMkZ/NgBMJ7PD7eVL6yIU2qjgBTw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h5kgqPrm/ghas5o50sQF7CkRrd0UW9+3Bgyf9II/ObYHKU5WTqvdQVx37RiV6Zuwx7jY8BKGUrC1
6GljDBL3LJhoaR694OorSigRqGQq9DlbWwvPpubN73/pUcAA/BmXyPJ11iAur9DDz8dL8u0AIVBZ
JMEcSp98XKgEOnXtjaU55MTSv0JNClbz/1GbpUB/la5GmUUPVd9VERL915SygcAxXa4efzVDfNQe
TDR9Cg+V+hNwUsZ4AL0NwCpeNAD+IBeM7wr73ySKSUjSInxlA30lGKpFr4nZ6c/01uzl+nrIAdot
iHHtG6uFhJXK84C4UUrX6PN4AXNBi1ScXRAvVg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qMPgyiJBLpyBHm6njnuRl+5NmZjHACVWOf0ME8HZlaAMEUuZ00geWO2DJ0BCcg6vVw2jNUSHe2YL
wAuBLQt46RfOun3ifJd0vZ0OhmxMdGpmaBkF+pDreoI/Y+6zbpN9NLfWQkPSbXW405FftA6mC0LY
RxeVKPNt7taRM3Dn7tk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GOYJBmvSniPrLCFEvUHh6c8XRUg3Opfv+CEOXcm6o+imohXua80ifxh90luGWez6hJmfSTaDELfP
EFF5QnNkriODMphgc0hRiy06hmsvCugkY/+lnM1+vmLXcLsYksCkRp1yvno838j5TK13b7OUrqjF
fpYN4rWrOt+Od0qedbEyjVw1DaVbqvMeSEy09YrquzpAB1Gn42zQnRqbZyB3P7UxKxd6Je78SneY
ZTMyCwaU8UpZ4qBnHHuRlhiw5mnZoM9BogaBHysLvo7BZaDOif/Zebq6qPrmHuj0Z7B8J4XLLpKP
kYrrZxtmMkKcHsR8kM8j5XlIL2/TVXXoecYL8g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QmPcEzlUpwA8HkI5E7k3BJ8/+g51Sr0bTjftiABHZ12feKb0yyUwc3DGo4XhaK2hwP9A/eEaRoma
DGsRKeLWw0e3ct2vRi8ep6WFdF7j/Iem/cY4NZlDwWOsU5p/5aUY6JIjthh9yRXtopvvMjCYzfsJ
/aV9biiKpCoceP7BX9BA/fsNJMkN6Uz53KSeUPzAHhAjmqbPrq1tftbyHQAdeTBIITSgKrbeoJwD
MluQlsoQv6FFc/AG8Xo3Jw0Xz2SIjACi5gXO0Om2I4nU923OlhwwBiwNqVm2ItyIp8VbqOkoT31n
b3utr1501a+m4vRbYf1P+coW4adHWojl7PGtnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 3616)
`protect data_block
iDYfqNwlpRopY+1YWynzvX88pK6zuDTIrvp/4Lrj/iKilTFUSYiYqhLUGBvHgum4P8PW6X/wKKKt
VLZyMOj+wQa540GH4pJy1FGqbGjpjSEpr18azZU2LoUTAdS56A51G9bTBop3+d7ke6H1HUcs4U6u
Y/Ki3Cro5pdYfVpAgEQhvlWJgTSy7JSC3htpWq5dVb8n5gYzweJSBOjt4aFYvebnifrkPGNcn1wE
WrQOqYYlGEhXRUmDtX0K6ea8tqFYC2SRRiYZM07QSmqHQVdJ0jWtU2ynfXi0ZqFNY5reCqNjUOUp
VPe41vaIQs146v98xYiM2YqOr0hnRpdrOVnEkSkWXRoaqjmo2G8Aq4AK41SsgBwN9VgczWppu3Ob
q/6IS0QFcCMQVt7gsN5eubMF/vedkdyTwjQxWJDdk8jFugbpBwnhuWHoYsLM+gzR+9Edbc20JIFW
1/a3iE5PTzXa82nOpvTmFpLMd73oqkN/g3vqg7l6cznKJ8Boe3Am5C+mzFtC4GgB+PE5eP83/q4k
PNKX29Wzj/Hu6F1e/HgabmVjJ8uRIUrnTJs4M59nF04qDyYoHUNp2UpRWD1LnSzEOA2f4GoUM2Aj
kM6rbyxGT/mwa/4VBquymxqogt+Z4jqWVdEa6QicMZdO+1UF6kjOlEkCIxtbVH7lcsQ5u7XRSc3y
euw1LHl/4+P1Q4XrLQT1rNJ7Wi7GG0L7SnCX0+S91G1bHs2pBs3rYidNdH9u/hf+RFFK6jx2h+Bb
egjt+FWDdEHoQ6BmD8ASRXrTH+p2wiw/3UQLTKCECXJb0QaqgtWY5HmEu3YFCIi1u13ROYLu0plP
RI1GTHZ7uzCs3exgSbU76rcuP46QwLbH2rvTuWu4UghNCCf/yxhNQ+Jv+kb+bpC/g1tYFUtUbDX7
xkeKsP1SA8zLWFj1ZwCo03QZ4AfYtw7skiE9lS8g34LtTsO18c6v0lrQtCZ9LTi6KeubNArOWwPV
F784iNftropHFoF8OngfZpN6xp3ISgCcjBwOZ8YyzEFQkpP5zAbYfVRV9fButzPR4x2lyJEWs8xU
MwQwOHb/9PiVTy3qKdPzFWvlPoyFjXS46i8KjMLh/0QtXJWkZtUOtVAbNJUzzQPrsE8Xnu8QE10N
VwsAdpSPCj8qe+iZfgVofo7oVoFp2YDHZ84aSY/Wo4TnjMWzgSP/wbYn4neDTls4wtsi/2TSoRjD
kD1juboQHfZ0GRFD/2XrUfeqSOW8LB32E3YWk5BWjm4SaayBU2tcWatxItMNjj3XzhXHdvgekz+D
fQeNGgLKFXD+pMJWLitCv0O7ZQN21ZKCPmS1qV7cQ2msv1TDK0sxU7/5dR6axzC9v/zsNahDCXll
j5Zz/X0DPSPbeJSN1KuDauHe+X3mIt9BZT+WvgTFVc4pOUSFXKXm7AkcsJ4Zo59ISDSio0j1BZlc
KhuIQntnF9EuSOcSFvUZxtks++oOM39shaVTNjQGYAy6AipIO94+5W6a0QuUSOOR+1SwaGq2rHQY
mN2HqnEqTMC/n9OnhMVVa/5vGuiu4N7yrA+tcMZAl7smegePb/GDNpY5SpIlhsPwA2waZFs7ZzcN
d5KYTI5vzi6bNyqjD9UKCLyEWgZgBMJYiIrvK8SWefYbOhdoXgs5SzGDOnJI+HWNc/GB6JyW9Uvn
8cIasL4e5J4q3yKc2T4sWh0KtS0TbCuL3LQrnlrNRQjBnFBZcPrQ6S+y1+KikbQRWddYZikQGU0v
CfiRYnJbmdbyM1XNKbWMhrWHFeA5SkC467azVqoJspNe0BOK4IhWwWop+liZN4dbZsb4ySYlvAtG
VfRtazKtrDBRIlID2o+69TML8tgadQ5IC1ZtVBcA03x3jFpe4q4jNyvGOcYndCDwakrLZqJSexOW
c7tcAooYKS8UzFByZo17s7j1wFw0kUqHcv2FHZlOW7EhNaw4DmxoppiBeWMO6oi+XvknjzpszV9D
lGPeMca8ei9AZKlZ2gnH9ntxTtuoyR/zm5lsHMNO3ZdxCpoKWLcO/eZzAmIhB5MWh/Q+SL8dCpAI
tMMl3N0XoEM90Jv/sdbK4OddjNvOmGkU0LsTEf2CmMziO6PkEjndYhPWSc+IzFxwAMfyE2m0TvJu
S1EI61LAp8eEtJqyK956iloxf6+tvyrCLMXA6MNCCaYeBNTOTDBXJOT8caG2uMrKyrBS1KISSPSV
tIYM9n8u65B5Wp7uJ8Jnqg95IrzSOCKe+ttrtrVfD+xlDd96Vx88qNLN397K3GfW9m0vTD7UaX8z
YEpUWnl4b4XQ5pPjtRrtGdufV6ejM2TvcRq+1JssQ5+7l7osszQ3GjPrOskeYk6Kfm4PVbckxNK1
igXypEpyespUdenhzb0OmNr7Hu2BlVd9rSvO4REhsKqeK22//2FmhQCUDrLrvh7B/8yV5vjJsweI
ojEhXrqJrnAqZ4f1puvWuQejWC/aiRIYllFmTI1CO+aOsQVWHw9dw0VpDNGeA8jT8QRQDSgX4I0L
RlpUPf/ztq/0GByQ9h9+4zCxj3EA5XXnHIjxEPF+w8RykdaJ0GOPOOmt3z+5QSUj3YDrCpbfNANl
qbF5J8r2aVqGckm7TRW1sAy0OBWFHplTgS5q2tewV1v3+0g+wvaSDB35/g5dzrT9m/SlqgoxJZyj
lH/naaoFI2NXP1+69ubwaeV92DGa1D5/gqFU7hSvTzbKzZTlrylYilgJ2ZqX87xPJUqbpMPMBNy+
PQjLRSXgzg5d3Kc8T58L7yIsDn4vicRwk99+VXqwrkCTmvzQuFF+dXfPCQgwhPLu6xiexk5CHwTu
yhA+bqJ8y7rK3aO1o4gfJEuDJsYzboar1cW4y5JJW6glx+UMVZF7YL6XcXKvd5yP92X5/3bA3lCn
fexli0LLImSqm6mzZcQv6frnXWvVnGZxf08u/w8ecKzn3WwRrqvLAjj4bT4ykc94Fj1FujUI2aql
GO0twZJVpL0iBBL4gR/WCZW5xU0ZOHLHLy27lmigv3zrOWbHHlri0QurigCIqoBDPDlSAIJu32ZW
OJ63XBHX1ILvfyOwpi5zBH9f01YU/0CcXWknYspbxBfjo1NHRTu+HVP+THCb487rF6soqw0zZ8qw
6ybcKUDOW19Z3ZKpPCbqHOVOkoVCP3Pdr7CAgzdBk9PMT5/98zcwNZmI86qv4+J/ZP2o/dFok2Uz
wbsnfh5gKnsSoSHEgF2NLKpmMcA50zPSik4FSmIThRycyzGrC4/3TLvw6mhkMuRN7jP5i1g/P862
M0O9VJS3MNUtlFmXpeQkCzZGhj/zYbR6r/uyhL7p6ThHbDTPR1hiAOz2UfuwcnSv9JNYiZtgLSci
dV7iy9hovvnc2Iv9nqtXyshIMxfW0CnVfm+H7J32YzbU8zK9JC/wppTwsV69SJ4Ynf+GJ4ZfZGhM
bn6MJAaKyQcvlPcL4Cfcfmfm7eHn6H9nEOm4UqAO0uw+4qc68v7tdw769CSyDVMwETfX+BZ74V44
F69PKuDSDxi5yql/rvc4/EHAOhClLhjxHTaedzUJmChMZw7F4bNdlWe12D7O91oaQJDnrSQbeLaF
42x6/Dzds5MEEtD1E/oz2XIez0xFU85mGsbvxUj5Ivy+aXcnXfR/Vu8kUjbCnMVzNG9Yz+0Lb2KL
FX+WNka8NoQIuwb7F100drtaOHAe/kVeMLLEgNnlhiZ2H1XABb/keqRT9xEi95IOBvaVL2Gszugt
Gkz6393tR030evjvEvHTzUwYZpopt34aNYbMpAtFXNUfMtVtro7q4SxtWo/5KcrlkoW6AEX6SBFi
cbx9JBjtAH4/Z0WCvC9KBVaaHh2Z8BKcKlybZVsauSVHWvyA6KSP1OXbnZLX9gYqvgS7vbnWP7Tp
I8gzw6hvovmLv46unz1TbSJhC2pbCrK9PTwm7pNH5kSEBSXHPpxI7anL9S/8jQuvZZ8re8DEI5Ay
N/dmouK67j5qbb37IW8UAQGl4Y8s+8qHHl3BHzqi0iiOSMBwPTSwKZlMmylaHdGOI0Df2xbruJ9t
4Ch2eHliFdlr1yxiAydR1EfrNibENA14e/1p3rJ+oeu7FLh9uNkbmxMJz2UZEYzQ7KAKPjJMN0qh
Xr9ESmhVYcNTLVX/Cuzu/mL5lZLHuY9Vs0XSJrtGOCYmeVD86LIjQhPNvCrZ8HJYDaCI/mPxztvv
42VK3d7ZW/EbvEHFVM9U909W3SisuCB6SvKwXSNovat6bx+KwcKjvs2sz22Aj/ofZ3dlhEB5WaMy
hgwJPOaaEG1uY6QbUkm3+0hPn7JtVGUXZliHRCQBTPizCRlkMXBdWW/xDzCPtYuzii7WuaOu/Xtz
rY2jHD8S18FxMadzb3e8fggKsxjtCxideYrHTNS0+YfUuOsVT4Gpp4Jy6DFxx6xqHpGAYJ8MrohP
oFhOdHu9uTTv1H9HSRCFUkZwOb7ErSi8SH6DvRpYsT2O3zVM6hsVpUd7DDgF3f4AbnPjyZnNSAbz
5ZmI3p55uJ+CwL1NonVW/LuWmmkorHEtaP9zoKgOYHWAqc/mo9MdpbyzkT44XZbY5bg3xNxuEzlo
5YrSni4hXsiAhICJLVViQuMkGXDSYCo0isEJstpBrSsUOuRkC7XHgltSi1/4/gw0TTDaQ9Qik+rX
1Nq88lzUEqfVa6ET2Lkn6aY/ve+/sNTaf4zBNZVY1AgkD5qE29bg/juDXH8Ckku4SUwfX24NEDF0
1iYt8GlMU7AIyBT9InaPRC3mA9CTkbk0nhrzjcob4OPSXzMQSvKaiWeFqIMHDO8JveRrXswHqUkN
CBQqVqPe/oDWiVKonLqU+hItzi1tqFYujg==
`protect end_protected
