`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2019.1"
`protect key_keyowner = "Cadence Design Systems.", key_keyname = "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hH+7Of7V0HrZN7akhr/PGWzFYMFZ/Rw1Y0MdJHcXbDfy25bCrbSAgiAHzjAOItzVH0GJHC0TwaAh
l8lQ6Djj5A==

`protect key_keyowner = "Synopsys", key_keyname = "SNPS-VCS-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
AmHoZR7VmEL3tVmWsOV6IVQew/VOu2KAm4f6KJfAzXGRTTxsXlPXI5eOmXy0OQc+dTQXlc4Nyebk
WOd+g7avEM/H0dDmrnyrAy4xkmGgWvy/yoSRg2NcrorlzU30DXGyLUL7cC0fGGT3+aYDfpalxOxG
vMlnYmB3ol3sAa02k/0=

`protect key_keyowner = "Aldec", key_keyname = "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
quTe40cgTFzwGZ4hh0czXTRPjRM65yQ2xuoMk4KWhGRBXqG0mDC0qybq0KDkzMvHMO9o13XXh86J
3lmXd5z2U8qbCCQTiQ5D5fs/vDyxOt2D8yzeP9Nz3v9pLob1z25U2A3IDkfdMys+0lSQ2Kic2K7X
M9l4gP8XjJ7XaZMV90LT+K3emy6GtwfHL1RmLLmz0wvq+4goCsSl98hEr1onaBQ9FjjXJSgHTEoZ
asLa6XQpuzHvUdrr7uow2fs6n/v6lPMa2QIEVAOBRHRZfcfQ8mCrRActebecw4kgaKOLxGzIWyFi
VJjLlE6Keg/yDxLLEGAzIe0fXmz5IeT0hi9g5Q==

`protect key_keyowner = "ATRENTA", key_keyname = "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
e0IXUCRiGRcDhitPNE5pcnOQjcFm6XyOGSyf5ehAs8DfcUjdAyC39hcyh7lelM2n1wk5DOyQUYdV
sH1HD1x890dqy0Bm+/WUTKfxQ5I0MfCdzTLMWpdnX0TYkOpM7Yw8f7rYC6qJM3409nB55jo5jbXs
BAEUxqIp85fdzNw1bsDtj4/QyVBwF3hP7nFhpQv+EKdvqv8Q0w3KT9MgfmK+tlzpA7nQq1DUqyYL
tY84oCcSfcuA/mVkkAZzSZD+v/Q3sdnagb4fc0bpcJT5TQnRzdluhqgGQtVo9Hv3B/rAkJ133atf
AhgpSKBM/HuMkZ/NgBMJ7PD7eVL6yIU2qjgBTw==

`protect key_keyowner = "Xilinx", key_keyname = "xilinxt_2019_02", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
h5kgqPrm/ghas5o50sQF7CkRrd0UW9+3Bgyf9II/ObYHKU5WTqvdQVx37RiV6Zuwx7jY8BKGUrC1
6GljDBL3LJhoaR694OorSigRqGQq9DlbWwvPpubN73/pUcAA/BmXyPJ11iAur9DDz8dL8u0AIVBZ
JMEcSp98XKgEOnXtjaU55MTSv0JNClbz/1GbpUB/la5GmUUPVd9VERL915SygcAxXa4efzVDfNQe
TDR9Cg+V+hNwUsZ4AL0NwCpeNAD+IBeM7wr73ySKSUjSInxlA30lGKpFr4nZ6c/01uzl+nrIAdot
iHHtG6uFhJXK84C4UUrX6PN4AXNBi1ScXRAvVg==

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VELOCE-RSA", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
qMPgyiJBLpyBHm6njnuRl+5NmZjHACVWOf0ME8HZlaAMEUuZ00geWO2DJ0BCcg6vVw2jNUSHe2YL
wAuBLQt46RfOun3ifJd0vZ0OhmxMdGpmaBkF+pDreoI/Y+6zbpN9NLfWQkPSbXW405FftA6mC0LY
RxeVKPNt7taRM3Dn7tk=

`protect key_keyowner = "Mentor Graphics Corporation", key_keyname = "MGC-VERIF-SIM-RSA-2", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
GOYJBmvSniPrLCFEvUHh6c8XRUg3Opfv+CEOXcm6o+imohXua80ifxh90luGWez6hJmfSTaDELfP
EFF5QnNkriODMphgc0hRiy06hmsvCugkY/+lnM1+vmLXcLsYksCkRp1yvno838j5TK13b7OUrqjF
fpYN4rWrOt+Od0qedbEyjVw1DaVbqvMeSEy09YrquzpAB1Gn42zQnRqbZyB3P7UxKxd6Je78SneY
ZTMyCwaU8UpZ4qBnHHuRlhiw5mnZoM9BogaBHysLvo7BZaDOif/Zebq6qPrmHuj0Z7B8J4XLLpKP
kYrrZxtmMkKcHsR8kM8j5XlIL2/TVXXoecYL8g==

`protect key_keyowner = "Real Intent", key_keyname = "RI-RSA-KEY-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
QmPcEzlUpwA8HkI5E7k3BJ8/+g51Sr0bTjftiABHZ12feKb0yyUwc3DGo4XhaK2hwP9A/eEaRoma
DGsRKeLWw0e3ct2vRi8ep6WFdF7j/Iem/cY4NZlDwWOsU5p/5aUY6JIjthh9yRXtopvvMjCYzfsJ
/aV9biiKpCoceP7BX9BA/fsNJMkN6Uz53KSeUPzAHhAjmqbPrq1tftbyHQAdeTBIITSgKrbeoJwD
MluQlsoQv6FFc/AG8Xo3Jw0Xz2SIjACi5gXO0Om2I4nU923OlhwwBiwNqVm2ItyIp8VbqOkoT31n
b3utr1501a+m4vRbYf1P+coW4adHWojl7PGtnQ==

`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 227296)
`protect data_block
iDYfqNwlpRopY+1YWynzvdDiz4ihvWKObGnB/CbpM0ndy3b8HYKHOYVxW73eYKS8P37UZXFbZaRn
OswUg1hlZrPhTv+I3noV7716GA6XzOsL1/Hbb8a/r+QSTiBjM1cm/s0KwaygyOzPi1DUt1mX5z/x
jEMKW9iLIi6aMkWTMu9VorFmWAlFyBxG0kAL83vGQn7sFnaAOfIoFXsbOcGYSDj5lrF84UJQ1Dco
SKxCbrG5B27bKX3AZ5Gz2/+NiAOSKCbfgNIyUJJLcGK4imeYkrDa3IU21fjr6KcBVqECNIUGx2AX
RAD1S9rRyB9azWtGqc/kMl4O1JwODzmv50M9WKHj0GBahn1ThNKQkGU/jYQ2+Bghk5UVGWYXxZBd
/LXmUcFPA26j2oO2tn1uivSQEtVWjMisa+s8E0MN2CmiqYSecIBNGy9nHaEssa9deoD9taggBszl
fEUFymtD5xN35b4q3rYEep/Sxnr2t8H+APm1f0+sW5laWgY3rLEHQFiFpAqO9mUFSMFCNf3ifduV
Scz3AquufJEmN7hLwpjgRQw0H3+pMOKxxx2mZf2uWwu/ItyREq+ADA7HOtnzHqH24xS01bxld1PE
YmoAwyC8anqztDxEIw+SyM3UwkmC/XT5XFtbBRK/JdWOtS56ItZ7i44mi9xNH9ulPqjDHIlHBhtg
ieARu8LUPlUCmHNPsS+X7X4D8ejlb7U9V8mFPi/rE4NtvGNyTbeOEcwjYsoY0nOqP4QgrvDt69PA
bUt5j0IKsOqo2vhqK4leGbrthMamcH/f9bJ8uivah+HtDIuy12Q0vQXjilNEKhXueDkeFqF2Q3h/
TEOcln6zJYE4tJQXpq+Xhr5Rp4sDPrivVoQd5+IaXoD8C486dYB8XUNpqnujdjWt5xdSh18AnrX9
bnM/vzcOgIXgK9INvqlYhn2PUOic5YOoJdOTGg5gWKmBsCF+x8mCukpSqiIotkayOuPfVe+CKz/x
9i25WZQZoqFsAf1JT388Nwy04l5znkF5n/bxMyJdatFRVmY0OIFscTzteK0IgS0WccSuz8oQWApj
pJHv9jjS05vHHKqXQ1T4j4vn+R0uAZ4tL4vV4sq8wgmDdwaWH62g5flhaokpgCdhlxcS6x474LGH
lTdZSuEbizGeLKtRV56SxG3RyeyWVEyE6M3ihlZD8fz4G+fVRNeXXLkOm0wsOISSyhlFPbBLnG5m
wM89Rs3tB5/2W/1Plune3cNM0IgVpdR6Y6cAvCgJ40LD4Y5nrdcRoOHobBlgGzKbwm5RlAxWpIC+
WPmq0SJ/Kg/Rn6Uk1b5/3m/i3KA5R4VTbXdfImos47RaRewrkVkabviC48ZDRdyezyISvTh3wmKh
9bStuo4CMgZ0LRwFK2gz/jnLvXkOTMA0vUtqKvIA9c2HQ2yX6RxFS5SbqCk05/QSc6r1rMPJX2pm
49IVQl5mNHLvYaTDn48kp6ug23PkFyz2KUAnxCFeitF2noLNGDXxJpY/XPIYKfv0KrBP4/cHIJNO
10IuK+oaFmaUebgRee3j+stv2RcBRmdFuXj6sqruw3WzcCM6dBX6szJtwHvPzj+IGDk3aBTXUiuc
YGvaEjbNEiiryIh9JD3zkIVTKKXx97Lf3jqM1de4gb2ALonh2pHBcgpGYIszqfqC5vQNaNECHAym
tZS2IEdJ2qsB4YyCLd1PQ85exOHSev029DaYJDuoj1KSsnIYlQ7nMqKGV+mBmsL+TY3hB9EZVr5S
vzfjwtNg9maT9mppDbgU8GoAJBZV2O7jUGxxrybKo5pDlxZZowahovASXMsYrQwzGorwNfyHsQs1
bJl0yoDlOG+CWmwLhITc0I7f2w9j9fLbExNA716/LrKw9m2bzGS8NKzBN9B0LD/AqbDMyZD5folh
DLr5ndCHRmQz5w01dI050QzGwRF4fU/FkoWqtrVjwMiKE6hTGwguaP7MixmBQ+AAvCMO1Hd4jdfg
PlJRzLDgXUX7Cz3HW42qQFIFBfWp+t3KnuzQkDI5qU1jVO2/xQwygLh6FmlKE40sFZ+Vh97Qtmhf
Isd22xLok2eLvyiRjosR4rVzc6T/ivReuSRIVQWGR/GTnJVhUwrr8fkojKLWe4XguyHeYcebNAc6
+7JvY5Kbyu++F5kwR3OmIDNjeVQfyJqyt1DMOjhr9aTVOZyHwhl9WTJShnDoR1vuNqcQPT90PnZR
9ljpi601vvuqtTrnD4oquIgJS6YJFGQRCXurVegUMLgd3lrYaTpiYFwxHqtogJugNDiP1c1Za7g/
VppGmy4DvFhkSEw7HktzmUHOFV28g0OqxE50+Syb8qsOmoFb9iw4Ig+0vHtbB24Sfi+wac/NRzuE
xn1nsV0W5N7UImPtuOpDPu6pmtoGJTVC7y7c7oDDgH0x7kq5yUlstCb0kTZQf2Weli3JR8pmp+em
jxhdoyWRTIgBBBI+lPp3ko3Si9belQLL9K3gZv0wrLEfXXEkMmcnCsKSPnJoTh6IVMZ1tQSRXJUs
F89shK0r8NT56BRm5C9g4vv6hypeWwCcY5hJH7UOzqdj1F8uH4EnhU9Md4RFqAi2BwCJ2vwFChOd
KLNl53AgHMcrMCXBLh87EXKY2EgJE+16KaVWpuy340+4RhbNtBINQ1L6oEH2VeZBTc1wMssitWNI
QtkqYwswOksaLEIstyYLFqsaPfGwZJLNnmQ+iCCZ3BwVWFJ7/ZPBAfW0bN58vNZ4QBC3sYJYPWcm
9nUk7YlJmGgF1lugG0KPLu+wHhyfa99yR1BNffLVxdpVjjIlW4F0G/BoMAyTpngDx7vJirAhHVAP
LAJX1Yhmekgrq5jJvFCYO9xGzTvqYBtnx+mP9hU1G1jvN1K8wyUrsLzLMQ2ptnGIKdempIIzbdcn
5/8jQ5/n6fTQ3flww/Bjrim6hJIsJOTm6oPcLky3wNXV20bPtIv7JhA7vTNQsDpllGBUEseIxawH
skNrbOCahPxb2YR5DOgBLlFbRRIf5HVpW1V9oZDSB3AvX+QYjTojRLyeSuSGRUWSxpz+mB1f8Fsd
M8a5kOyE4LYLYIU5Lbd8UoBXKSm60kapwkkMvNg1pOBSfMp1ino+fSL2KhR1PX8Qd5xKKwDPZXCu
wPoIt8zCq5khK92LXAxhbuVYJvkrzwykg6lsIzwEDyc+dClGpVTifYzJgoXN6ijy33wRo9NeR5Is
SB0IMJigD9JWyBSVM8AUnRh/KuhWk7ikw435a+PiAiLok2cYFkOc34bZ5OtoDUL9gcTufPheCKKc
YUOuxv4OqKkPblMnh2aQPIVuAW9PfikT06gf+HtyNRWwukS3CPXK/Vv8b6hlMC9AP5EhzHkugpz+
8vwh3IJDhHYuR2mhluD2iH44UshOWZl+BzFrkmUgMk3sx1z/RxgtZ3fAgNT5SQKnlbgYBF04tkH1
+kTi5XRtU3uBJmlhvqSy8LcP2euxd5E1UGhUP1cdLOXvedqoC/lNodQiSBuzBXdAUaMZuo17bpgN
TdU2++jHN7SLmIQKKxskszfRycAmh6w39Y1c4HGNrBufnqSxgiS1LjeFLuKEF9ZJzea9tTH/AtlD
mRJSLNFS6tXDV7dN0MsoV+xKw53uhlG7YOQUP6RbXrdhbGUxy0HKuhDRjRny+caivPJScR+dcyq7
G5LlcCFc3II3IUirMwnU+GuY4i5HGFAMdSEgebATfG7ohP8rMXQoC5IwJIgs038aqBSoMjJmWUYV
8w2GrK706HZv2VkKPeyt1D+VGuA3g3ilKFQ1NoWFeQ58n49AbUvK+dveuSZzc62xaZreaeQ/Rn9F
mfeW7+YapXOBniwgiIXUFgX5dIbIpv8aGGIjKC9wrvRg3rGkpTPyHlRm458Ycvg0Z/qUuCsRWf3/
9r4m/aclqkcbTDCjKAroEoc6VJ8BGNuo9t93ysStOX9YV2IBU4b14koKN4J+jr2yiEXvzQUsjOEb
eL/8XjO1wwxDhzIae1q0NJTm0ndxsu2E2A0+uw0ESuln19fPx9sFgVJ9fJrnWs5bXnhw9SVVAfQG
zEUwMtBk1VTG8UdVClfxKbLheG3smBKlhMqudUrlM0XelP4sG8exKSqSNmugXKnYuVQCi6oUHI2F
dvkPgiD+97tSVE+xZeRsbCrNeB2+GVVHj+DntY65DKfRTTnMeEFIZOoRpZzsEeke+WFHeH62xM6a
w8YFjBiSKHyJyswB+1W4ASuIHJmRIpdwSwr6R1PCT5FxDFbgAroTstH6+vE9jMfnSNLWDSNRivI9
zsXBfGlilJXqkchBIIWq+ZcY30owQVArQfbMmEEtvawjfAo4X6rldDRTqS6bTH5NMnECIRCnavi/
/osIplozlT51pFcmNWMbED83OAIHSRqKhV/PqhnLwZdvQ1fAiDP4N/1wyoXaUSBYGTaBKKuTgKZ1
SA4GzaRueeAoFCSYbjD6JJoSK1MT22Q8M2LsXOSBXdgehAuiCvtFa2OLLCX5I/97zn1MhcuWf7zy
3dTnT0Z4dp9LOO6VEqnBRjc+Krs/dvY7LYyySMo3TdzFOYYxnX5Owkr+sA1T0t38CTM1yqjTqiCU
vZFhLkmK7fs2BOQVjsAfVvj42toUmXRuQP+ReSUHXK8F0pVRI73M65G+BojTwBWX3QYCrVQfFLe3
6YB6AXZRDKuup+JONVRrhSPBqvOVZYR6LX9m0zRrScyi4QltNg19chsB4YSK3qdaxRAQC4b9L8df
PdOEaVjEAEEuAeeuhGDy51HZh2c0W1xSjQS8mxnhceOGYBYPEdru81bkmI5NJYTuosxU1QzHliFJ
aYge/WG3AYW0RmIBfzj2Hv/cL8cy6yytnLRdZ1NlY1J2dFNEn5UDgNZWxxj3CIjLubsSKPT+Ug8q
z2cxHZapcE67rqmTqlODyl4KshXqoOb9orX1gMJZqT5GfzwumRA8mCviujN/0cYM2lQkPEB1Ia+X
TNXzGUFx2Bxw3i0aoTomrI9ACHPEX4oABjv1BhOGrQQKLmaiNtxe/AXMJ/Z/wBnUzkFa1S59GJTg
DBkWfH5IU+NntOS4nMDiORcGwVp5FCHRTwIbp9dNUrvCFqUDOfOizjrCyZyz39eEBfxT1Tb7h92p
PT9vlNVcDAa9LonZl3ie6UmFqhGSfclEjIr/sjwg0iHaX4Tca26H9owr5SOEoTkfvbXfbBNeFWMV
baXk9tGqY//ZuaKX74jLzh8bUjBP3TwA1oZMe7ICODm9e884GdIWEj+KMgMbmevS+fpBvR7l3Qzl
9flTQ34LU2Lu7r1nDkGDcfh5eHiby6zYBGkHq2tJeqUzhUAqj5pAwGTdQdUWWoee+cYDvT/jMIDQ
YVTI2VepofbM9yVCGBtLqC6cPIujwkDsctCvPNMWIofqcVsHqTlUss1lKvviZPml+QW6fc0TFDOo
RVBwEmPTJPloK+x+99ylB9f/+IOpf5N1dL/7sTzslhUsQu7760yA9a/wabQO87kdBBs6OavVRh/d
SRTz7Est7GWbjhKJvYGfj5X133HptsXR6Fmx18TfqhPAi6YUXkIt6gFcyMyM55yuImaOpp3rs4sl
E8iXxrMQGINyqqq2VCzXfQxWnUQTYWBVTOIbv2LrBj/ulmryndXhAC20UnBkdTW8LasCmarErDPV
1j+01JLXUkPyaLc+JSC2IFnTi+xpc1qQJ1BGPan0Tdg4AtwvJTUAs93kPOTZND+2paMpD6IoUWTT
m/OLXfeh+JD4pWOXNpgzcF1MCdP3Al2BNkAYBxBDqsQgTRLCC8AKcRwlWZjDbnheWbAlMe9ej6L7
Bu3TW3TmrQv1aitEZzN5Z9IsWaSvb+PNxmHNMgrAuo680sN4uMy1QfBIB/KQ6h2sfZboN5/CT30M
8Upf0LjHgB2HSy22yPbqCGldwkyKzO+jVloetgMA4RRiLxGp/6Wzfe2NgIIm8D9yRk35nAHlqDCq
7ouLvw3A4CJKdMFBj7V+bBeztyOKcZ7HZnnRBknUoUPSCKxfbhqfIrGe9OrC8XTLWs49sZm6WnzG
1VAqKAAChbA7skjDbIwqIDte1ThK2rn9Xk0xXTrosb1WVRHJ2s1x+gCe+WM+wYg/7Gz0JhaCoDJc
3+YNOfNVwuNMmpp2HybWk387h8xdW1BzlVnFp6YQ5EzeRYRhLD0mEhQwVY9vkG2A2Oxo7K3LbzPn
2zGdsQ4u08nnPM15xzTnfXANdAo3fcWg9qynoos6jfWF5Xyczv6rq8era/C74xIdnLbyNLVIC7zi
wi6JkLVwQeuzlRbkAA3TdR9rso7xtomVyYNLfr4jN/0cWcpkpRrj/wTfh/vDffeVAVvK5JFaBEvn
bO+vtJDkgqLaBEX838e5C1aILShEg0xZ6SPNZ7UrvhAeZkb1gVAy42KeuUs7tt8OK4/XiajHi01U
sCCfqDEYCKxyUImF5AbggxLx9lESJIHRlAaBYxHWvUCJBPX06PmMgc+Ognt/dOQVxmIMCuKMzAkD
v49DHdGwYVc7WonIWPFkmGEKKjRBFSgOsRP9sxwsjcFMz1CZnVCJcnrNkTCM0cJUhJFwEe8Q0eWe
o5AwPhsIwEVWyba8n1BJdoEP+7ZnWkxvRPk3eIsAPnSxeVxxJuKebVvspeQgQq3cE2jTOPcvhLKP
4axQy5w8t2h4AZ+ub3Jt/oAxqQIJ4bGNlR40k9t0OxvfkQKptXtaGMAuwBANoGElc/oIjieEE+a1
M5BTBFkUZfqgcamJladEYGb9cvFRJCb3PjlgNGaqIQ1gHzYejaGeb4ekWMbYW1vpc3Dg6lFkuaKd
X9B8vSh+Z9wM49bFLITisI1QzHBYs6bNyU1i59sEk9HGioDLTqhQtx9uJwADu0TJdJvY9gruJoZP
ptD5baUriiZkMSe0i/IobjlOi6dW8GqxedCb+VcVjFHMpcWSNvOws89/EXd6EsoF/kQcQ2ljq4hl
fA32QVDUPz0Bc8uXH7xQnZoUo6aJODGPTfaJ2x5sKGSoYF57Q9qLKtuulUG0xgtzDXJTNqo9yyrR
6KNDVe5wgIqOAeNtsMeCmipeseL39ZHGeRI2ISHgEJbNV2afL/yBAQr034/ktHi8/esVmsXfrlxy
PejgORUhDFTMjDyOlHBGs2COMGnwldDJTvPGAKW9yhHSR7HCc2f4Zy5u1gB0ETJi6D4rAxyBhWds
iX+pmek2HXP+FbKN8kgDFoE+KLb3R7fxeXbzRdY+jOtOcCQa7Fskqt5jzojv4gsO8pb+oWwtWcN4
KQBM4zQi4hnQsXVgEEknW6FTivogq0UB+2jCWUnsnH2EtrCvVK15K/67GfIVb9vlB8a96QJxxAfN
QqZNtBcnviLrhRRRRgrevRxHXeFGrWAAjhCNKh5qca2vsOWIrYvEcfJcETcaNZpAo2XELMfNRbc8
Fqr6rwYQlfyI1Oy5Skj1NYj4lCFgYosdbOJg9OkGzv3w3GosR8zUc2j32/IBFE1pkSi+6g2aJQjZ
kHDYnDgkSlklvxM9/e1u8HuJQg5M+YFvDqrbxJrSX7X4OK0AzXFWyV0FKwLu9fJy/5nc8QaTCU86
MtEnCXplaNBGZNJiFlZuChkn5dEJu7Le5USsvSrL/W4aGA+I/hS27WiXAXySW3exq5BreAfZLBKh
PomDqHg42qNc5ObUg9bSCq7u1HaHQoWmjdOzjKivgz9OrwKQ6TXoCxWPB567Ni5SRC6BlNuo2fDJ
2QJX5oCoKVyeD3Jws7t5N8Njw6IhsPg0qfaYyym3+rLh9FNUG2bawHSvrTBHj+xqA2RQb3dxJo2F
YQRSBOBe/r22fi05R9hNZgmWyw2PInJWc4D8XZCq9iLBpEpMlBracPMHL2UvJAGXKtRqHqD6wfC+
0m92WgB8t8hB1ysK+2HZyaK6vnnx/FkRAeMsGdCugddz8mV+/eSkTCSUWS+BgMxVNP24U1We+3T0
V0n3WEhwpKIONKFkmmgD682Cs8r/32KfSb3xJ/VsHxLDmIhWVQwVYPrASmnqLIjzpUdUl5mY7vN4
sZWc+SPp1grToEg4svFgaA9N33VZBkVigRGlDa++gramQn7Yw4gLC1d3LTydmEXBL+gvsRWDOzLh
PFTNVnTqEjc+n34XBdQvjGBkKnGziYBcEOZKKPjdTiHlsjrz3rri2FWejDn9wQSTgVk5OCEOcuk1
KA6/a7th3RQgieQveqzF4lwGjk/MoK5wUPEcRYfKD7pvRkK47AlQU+vsfPsu3KDsR0L9ZiXKLMwy
HDGhiff5/geJB4HWmz3u/EvIdjz/s3bluCgcf3KwDRh4/Z3bf4lZYzrcWtjfjOvuU683OPFmOf2m
1NMXOIhYV4zhUb88M9oMzvr4AyvIA9HJAj0wI+XjPZXSsMVM6jTRLNbem8T7e0ly4TV1OcvkVJDA
gOED4nGzgNFZ1H96YwIvt4zfvCqD/JA57cAg6b2Vts9Uj4ZxofHznt6de/4/xVmrmbl4+n9Hqs9o
Y0tDW5KTPjWeY/CJ20xagwrwv/PEQaTFtbhxylKQAsXbEsvI2DKr9nvtEqqn1F3Hn4YGl0qkZuck
ZpiNbohia5nr6/NAQ5p4Y06UsVplXLTCOIBY4teRpug5HGbtpI7pXRF17jRTUN+R9hSulKcQQwJM
kX9dTtWY0atGq6ApjZ6UvDK7bXlHw0gpKWDvPfFSmSrwPIwEeMH2U5m7hbn/6utJCOTC6LBrVWXr
1faMHL/W+kJBH0faOh+TSo77W82BpG6skcEzHj+FjAZcLXLXHenGhQvg7lxvunklBajj19ARAn1w
wcex+SBzk2uDR4V5JvoT2V9QtE7Wq/8osMibtyAdtJopQEpZgtv2Ikls3yFbbeoF7XCEzDzcBc11
/eS5Bt87sobKc8Zl9aD7n2E6ee/i/hKhA6k3ly3VtrXq+LG1SS8b8I2kCG/v8pB8toq544iHmq7+
h0lI1mqKHn12nNM4AjZWc6MHoQkcxy6zXIUndK3RNWhdoVKTgpM4Me1YFGQmoNVNOHYDxzIQ5uky
Eb4zyykHy/0ayOsennAoVbtaKGWfbS64eSWkhv4bqVl6qMsADz0xDsSFhTeiwqNYPfJu+gvLhcW7
12xOrTMd+7J3oPYH+ZtDwZ4Ytp3fWP0t6D3o5zRsZsxm4ns3PIg6h1GSrQG5wnnhuQqvRFfrWPy0
owciSymEKoF+ifDnTLSl4Fv64uJYSFssaeqdWcpvhI/22MBq7AfoQgXFKmwrG3y7q5rFR5f1dDHk
8X1eHsCAOeO0/Kr8rD+1HBs0hBAYfOrFV6zWRplsalU3N8wV8oCNFNuYt8gIOv9B5n50uXVB+7xW
ZBClD4ukVzeGwfdbHHdNmz9B4dIIEATY9oE3HOmNgEyswwJ/LGULPh+gyRyq5I/9F3/G37Yzm80F
o86NZDFIMRWhyWFEHS8rVNUuOh0+wyEssspDbB27EaaVUrQz96A78pKA/9Ze0iewYKUCf+OZkHZq
yL08gyFFDUSHYHgt/T5TCo6nM6tBUs8cO0OiREws4Zp3cJsQkSorw/YDK8r9sJejin2z10Ml0I/h
ecJUfmbZvoiAVZKmJPmbmQI+mUL7NfKATKFaBfv1BOn8ps6jXi27QBx/Fk9grzpJY+bT/CLv0DhJ
eA4ejZ7X7CFTvuamyY4gQOzHGSwATuEG3Mb1wUnw2rAkaNuoF2LBYsN1IP4yMQoA6iHpZBR0K+zM
obt3hBoW4SCxTjjRHnS2PAqCwbM+42nu5zcFsuv7XGx82Ky0w98d6RuaTEggD1JWq718OnhdvY4Q
UXM/9UIteZWHuwwckNstvBN1AoNEl06h10fuvSq5z9NzIC/kUIxvXJXJGq0YDgMnzEYQUkzHF/q7
wyGnQOgKBAiSQNHqQti5vaueXsLa0Ai/gcou+MfoMu1yjErTC545kWITXJ33VTtaUoCKaBMbKcu7
C0Lz3BG+tNgm+b8TBAyoSZWWDpkcAkyq52SWJw3dJ/y/uykhJGKRuPTz9Wf7/nFuCcmSOmQrO7er
PFlqhwTFmgLW1wgi05/5M8jHeTAubbp8dXfZDTM4Dkb/eWYdheWygWUNxpICd69UsXD5Yj+xbjlP
ekcxlOuJJkt3V/B4s9Ef6DLYgxYB3xKLbsgKSPG9aVTv9pNfoigJIjnWeTtv9/MLD4R3lm5bNUG8
CdXHGtb72mxIMmhTmA1Ygwoxpy3Qa8kJnXpfqI0RcBOBVELZ22IUuNEtZNS5ZIvTZlmW83LcdZu4
qn6Dv6jdvlgb5lvXttPWXfzLBKmmsvUWogAUgCNqzyqa8M0EWsJ0rhyZMR8hTvxeCIfnGwqJkbkR
pZTPZJzpEO8bFEY4Rfx0vCL65B+oOBItaKRnqcLGut7t5omg2NdWJLeaMGl7DidPnOETSaOHrygy
sb7Oc00fTIhHAE94elYtElscqidb4Gt2bSdSwwFK7+TB0Icax6rZstfTVJ0l0+3kOlg7nfUft0pi
M5DpvEu84pvWyMkMWfWFz1BvzQ9HkhLqgB9N8shkHM2NdgJEE00XjHQo5YeJa/M1wUPIia185h8Z
9lMcaAvYPCEMIw7GkgahM3sy1v7uEApXJhdsNJuxeLrgKhVSdY4Tgo26/zu7r+p5zTY3tAMj4NPG
DUJ+sNjQlTYuj/0fLGd66Y79k7lYFlz0ksBvgfFqxp9sWM6gOHxv3cWScnob/88Gyv+poVQTaUMp
JI6xJ0xCbIi4oEu2JqgNNaWFwmCvVYC28wGFcav6+sE4nGGpDQSMQKH2Xg5zY+WbnZEF8rKcLbku
0cXtdeWLUskEgJJG2InIcDhS++qVHQefbiuBNYXL9eU9cnEM4XKEvssedbeFWsFiH+B+yGN96dYc
6FG+E8lDvPCjFSEbpYfkRW38EWI2iVkElgU1yu8J8KViMl4itEWzMgmqpUGR3vG80HaUpI3EQN+G
o7CztYVatu8HW/VvysbpF81UTTF9dYIadmwYmKn3iu2Z014lkpxw9OHe5WkD2BEHFE/5usQNMQj3
9hINqmQ6VueV2fXRdOdfD9547v8/neBF2ljuO76eYNTCAA2irnWMjfOfXQPBcTNDXIi3Hx5LiD70
8evHWAFm7pwydEgTS3MbNDPhpeSJXNhMTOKHtmNF/hE05bMMln9SHDHqwafNdvMNrphcpeC202k2
jqGYPCEF8dk4+az/zfJY/fPxRotwKYMAvYJ4W2CqcX45ky2eS1Ap9mZcnGFFMdMhemTbNO4dhizi
2bm6AtYoROPVn0kCHSGO/1+47tmIx21j8OaL+m3z3ddFYkiwpwW2rOaow7HmRZSLw9weGGp8jaGV
HPPm924uvzhEQhlsBnABNOrrIK3wAZD99nUz8GvrialpJjKCN2EwQUI7LtR8/urY7ffX5MP/yuCn
QmIp5nQQL5tCdSa1nVPx4gdwyuqWlH0CRIJrgs+zkjRICctuhqf5wwAkShjtzDqmg3LKVhYSDwoI
sW/SM2YLiMmqpkMZWoW1oEw9yps8UDXhy1Ow2EirBP8Bn+qDVBgLUWA6xSKc81ZjsNLvMfhz76w1
MnaUlHAfRo4uOqpGs2VWq/3laMyXKwdgeSPKhahkrd3ynqisAXC0E42k5iO2D5edzXsSdfvBHziG
uKPdNEm7oungJ/XzX2Ex3SxAQbj37h8JwLNDx1Sjk13eJN70TFwCDNmU5bp+jW4HgNth5AcNBvYs
31TZm2ma2pIwPOwNPnMgVoR0pqxYIFmPBPmRW1tM74BDPhd82QMaNKnR+kjyNhiJYPuFv6w76a+7
lswnL65WVUuZIhTq4Bo12mWulpNigputkp7gze64RNrIG7Twr0KXuAmQ2neyvZeJ+vxkzfX6yhEz
cd00VDqxmPFTlSriysrOx1PiVstBsXQA8GIRDOSjIhz27ukrIkZw4zPXh0xAOb09TAp3yIhKa6WY
mmsI2WPH4SHBP0D6D7HthQdaLmfT8WU9vJwzgH+POdCWhAtLe51hY0bFVfhExCyydgmWTNhB2geT
9wtr5G3NEvVkq/5tteZOknowLq/NcpAt6JCY32Y0AxN9sxw9xlOm0geFx0pP+h9eMh/wOMXzI4/D
LLyZ1baPpZFZmcREuYCuQnKfkTD2bCttJZ4KFoIcHZY6jGgn8PeuBUGSf10q1LTMAtGQ49ldAwOE
mrlkJM0Y9soJMr8CzlX0xEFvEnvHeM37KiMotu5vN7kaYxT/5WtBljWYGCm0lBn+Cgm0OidC4V0U
kF+743626CVbKXo5i1crwerG1zgD/cPdh+AxDUXMwPS0UrGpSak5vvNZNdpQmS0ziARyKOc/wSTP
/QXwCkZ1gZ42BGonHKqf6NOrPFaHAbJYHQCotVsoFSqWLbp6QFKDijj6ZoXldy9AhApPA8ldZyVk
8JaFP7sl3Mda+WlJ2KCCyP4YR1eMlQl/oMx8ToKIIhUeAzskNudIaoFQRkGNz62Iv9qaNPcudm7h
lJpiUqCtS/lnzVQ0ZhStt7yvltG+gIKkqsKMzFxn0l8AZSSPNebzjmjRtDSijnW2NjUQtnz3beGa
jM0eqa+q+0OJojLVWmJzQtr/a4ahEGoElW7vqvyPqFCK7wSRyyE/TwK5UH2oMCCksBPPHRoC0c5/
FMHUIJ5zLLkQHJjwX/9DP0veLnEIuVlHESgKOtVjMZgQu4dWlpzwfnVJiw8yN9kmfvkspeAzvlDS
S6Zu+3v+0ScgSYsAk2IpfTlH/KQQDJZpKIFeRww2T9mwyvL3KW70KIaP4c7OmICiZB0Kv1QVdGFo
IlQD+lCZ0XEbZSxceSNdqzZk97Wuke9w/U9bRk6mrcRtXI0k6ejeQEXJP4MW5bZ69hp9a8QKK2ek
ZuhNOcXuirfilBJ5Gz9rYIwD2+75K2n5s8fSdspG9/VtqZ9dBqImD3vWg5nd2+p1dQ3ed3Nbt95+
Nw2Kf864dzEZHUIpgQFIHKATcJAP+wwuBTq9HpoJsI/hROZaTxT14bgdN/slvWjeG6nLtCJA1plB
ZLZKtrpbcTydeU3Ns5vH0YAjNAikfqjVIoPIr4ZsSkY5JgN0xcRoWSnC3W9VcbbGNr/0gUEXyVq5
VNZMVTXc91zYHOLrz89NvLkHfUgOried3pUYvxSFGA7Yxk9g8xCt2ptrVLBe7dhCDNXT+u+W5jYc
qqQLjRrOaiLoKdiPzIpkYZDHAWKDAcLtZAyR+z1xtpHrdrEpUrH/3sHzXtxY5BenoucCoIcnUZGl
GC2/+Kwx0gJNF/jMC9iERLwR4J5WKreHGYHw7WRdiSQtJI9w77ufdUFDgB4ZLFWDbRyizC1SkROk
RPI5gBvi68GQB1lBvUDecydEB1Q643Zijq0i4MVT75H4G/ym7p+AMicIA4xvXqh9WUP7QhFXJI+A
Lf1JHH2HhnIoOWEji9JzfgP6opCk8RbMQUbQcu/2EmbMW2JOnwu38r3E011L4mg47pHWqwfoytB8
rYfkLO+YKeBwN8wsIJSavYPy5LNpWJJ1KL8rMYHrfh8bpbkZt840IXDfqpxeK3JxC3R1T4NDCtko
RW+zaciLeT1na7nB7EL9TrNHUpgKcDajW1GTRDREn/+T5vfVJbbtNcUCG6EybYDASg4P8KBdkQxB
JEAxvdg02d8TT6wAXsjFHpcXf3M2LDfk0Ot58cD+ikwKnTz75HewPaf4FpAYuC6leppi84tJ7nJF
SFMwgKSNlFL9xZk3+k7rgn22mhwAIk2wTIv4/6kEPlPSMo+y7Vfpc2fUJlIAsULNfaX4eg2LWcnE
RR6yrCulp+VSoK2tOuBY5Jb5HYXRPhzNLPAOBGo/VDgXNnKG89IJFYEVWhX/bmSWtOB0106lt6Ht
e10pEfusp7SqF/Pwh8cWA5man0t98E6RmhXFW2qA+vSGkVXBqJK5MhGbmb7XSxQIbbfWd8gbVmvy
5eZJue2jGDupv6F8WVbi2LJdmaDReATYmyf1VvWLKzpsLSPF00ErSE3Anxn4wwYsHNl2NKxyO2VE
Pl1Vw/HOT946fxyp9iZ9F9Rs35m8YIss9yVAOYJMnzt8hglViEitqvmjbNBxBvv8aRiNR/K0Mth+
Yw0OiR65RZZFwBt1xLAVhNxlr0b+pbXFskdr3G8VMXsXgool70OleRLuh9tMKWU1xSzSWnrKP+lF
g7g9AlwGYS5CncO5k02GGKECJ8Hzvr4p83Q1J71hL/cApg7jmYbZPwNQ8o8DuBtorN/lJx8FEPQM
PBjG7a3VwVyNYSSsy8tVeOkJT1Zr5F08HanXYNoNkiqqfzqZQLHN6KvFMA+sUHnVzD+yk2YBFeHX
zjpReCIoDKlyjlN6al5dLZV4T510kkhpnUBMSiRMvthhzcj6GaoV6BrCKPT9iUAunwbIcze/Svv0
AwUDjyLMGQz38vhxJ6o+2/WZOGcGNpBzmUprmjFbf06AzoHRlp//P97bLzD4Aeq+sNb5P4iLv5/Z
Gr8QrPdIJl/UjPx09NJZ9AwNv1NXatmS4ZWYI6qKpPTLlx764Q3D+jMZ+p6CDcA7LqiWu24ZmpKt
eLIdgHx6Eecp7TvllboqFBR2XN/tnH3NRPYVG0p1wsQoituk9nDeamz4G8k+Tf/F+XnP0koInZJk
/8CjonREcuXh6HWvEt38VD6eJl+nz74/S/5GMJ2h3RbmiJys1/2UVl7rrF/CRjVT8+79FzkbQlnE
rEi74dOTapRFbuHlzOg+PCpUG/yS1ysj4fAKW7HNm1ZuVR44RsnvDINfBLC53nCB1myLHGttPoDf
p4HMzGWc89em9GrfpiMgRIaPM1Zedg1aDT4HkUe4OmeS87e/ByKj2C+dCr4VzePti1CTIQ4PpqHN
LLJY+h7kxeRl+h0jHOYjfSoQF8OLqAwgGMjtmqe3VmA2JfahYCfp+98okwCGrKszFNxxOtXYAsv+
rBDe0nkCGVSnsnn4TwlIsjXtFabedROoXLtzyBZAwcf4dtdJldwB07Y3cWil+XTNf8uF14s+KJ9A
ef2XoicJxcuVe9Hbx0bV+1hcwO8RDL8WP0ceyHKeiXXjCY03VGFxQgRI2Y1+dcfOXmieolTJhyZ4
ss+uwSykuIQEd3Ary92yUkPgSghX+LfPrmpT7PTeF4VXGfKiZySEY9YtK9/WakH40fAJOcrZq4lB
XLhbJ7wPK10CnX0NlhtRLTycybfoshnyVuekYRcNdEKcbR022RxsXrq/YHnnDNV7fCgO4Edf3yhU
pvYicxN8mxL1ABLKc1alMj21BKBMxiF7CqtZgc96sj0pQluGHIv3lpvfhHIBi+M4GsfLgdJXQNnN
3/fWBHz5XPl9xYykXnzw1bWNKAdeUk4xKjbYRyrmnqwY8a6mvks8cvnBVh8oITXzyyDWih3wpB+9
xu3/fdO+cYN2OJ4kJ1jEzj0Wyztl9FUBdrFfv4gTbwoyrRjZrbiArb06c8i6lcellS7ZJP0D4smP
Rvy6Kh84CdPgD6t+bWW6nE4IpEgMyS107ufOthqZh/+gXMjO37HxuCx4Be6MqVYCwxNrs0j3Saph
iIl3xRL5hI4kDcSVhLFH15ZA1o+NjjEu44bh/uceEZ+XtnuNsvNiJ3LqwHhYGOuYZZasLh9XtezI
lSK4TqLIrCosvfxoJgLEQM5dj24FQ3LODOotwHIF/kGO53sbS0KkTecpj6M2FSTol3nOz7CQztmG
0a6bYRgxSMfTxu/4NG3QYR96M0ynXXK8ESkCBHgNrflLZf/+EgDZh066HMTa/Tx837Rila19ytAZ
T2702QKlFCpW39dsIl/dmTbuesj1tol1/TFtrmKJRt8TWY753S0fzKZA1yeeocQRsLs+Vx3ZYvNU
VK8t61SFBtiDbGVPp6x15XOwyEtrF4682jQrkrd74xlAPjIn9tKf5tdZ8RmCF51zgqPi023WuAGJ
DZ+hf/ILpbZkCOrmg9laWb1PNIDJJ79JFS9WCQtIC3H/4IKu/HtIQ96KYfI4jOTkPhxsGRm8UC7C
aFvobCxYDPrgm+Ls2driAo0jcd074hMtIuuPbrFxmUP5WgPg0KYBIxEg32LE946cM/IHdOxgGcO0
rrCnBEDXO+jsHppa1Z7kETsbhrgpA1pGZQ6JsLOq5lM32XJs7GxXeWKRa2UAyrTC0dMqMm7uLeMp
iuKxTtr0pzkQ8k4CAKeLyQigVAdzRpW5XuFjHK58TunMr3BtG9Ij8Q8IT/G2YDB74jJdUWCVQhwT
zsJn196Bxeggs5w4r9fSkYTk4qlDW43g2HbRPaxr7yc7o4zuS4Ps3BaWQR0FLbV3OWfy4vA9z413
IdP6/erPI8YEBzQurUsLkAbnSRUctyskn9aA512dUlvzrrHzoW0cLCC4DJfujZasnPMDOK4f4eob
+VP95t4efqtfHkdEG8HFltjBp62THWrxPG2hVX4mxASxGfp8DvCgg0wqaPoV09kqi0dy21MbFbjJ
VP9NYyXafafPQfSrnJYhQ16k9ygTpmZvbE+HJ1z8y3FuiBOOOnEcAA5UvsXiQnbcJhLTUVClP9DR
WhJE5EcIlaf0XAyK2a/F0wvMVjA+rIxT5aKZ+Yn2FGqp1b0TtJ8Z1xrkMuJXkFhBaYltKVAsCQnf
9gScEjaXo4/nK/KL3vX5SA8zIpbKfCBFknu+rZovqGZCo/hLunLc1//tNkr9WLtm3eR26/YflyF9
b1fw2OqJUol1k/xGfwKyvfyCi4aVwKfYXhwVw3TkuUXoonb3ZrSZShdgKOAcEb5nq6yDiWQfJiZ7
kkb158unVatr+npQfoary5AWs64TKsm1IST14G8p8QbvBCHDaWZnQ+oXjmKBlLKKKyYHieswoNzq
y0WLVuxHD19mgNHma4x4+a2FiSPXabvA1fDIoXDKcJSZewgrgzN3H5hgwer6iWU0r/WdZPeq5VhO
wJsjKplNhgMFCS4I+fWelCRRGPMHD/apT/OoNXOqm+El375JCu6gBUHSnrcUib65v02Ca8XQAfOe
cHSQhQoKQrBQ5mEX70of1noSMX8p+3KfDF2KCwoOepGvox46xpzCiWB61jquhyZ5gZYUe6rC/tQt
FbW/PkoQJJk9kiuybxxIDUgyZ+H1iWCJf1ClfNFGUOXIYkAthplRzLuKwtqtin/4HzXUiYhd3MdK
RmMTQ5nR+Cmw9Tpsnl9tVQQbBahH6AgZtn3s1ziftRFIENnZqBmiXzZ3bCUwYUhcDR19h+xf6hU+
0skC+PlkqgVd4v0/wFJ/mEEdfTq/9PYjmi+KeXOKJyOF+DyzThDXGFu7epvjr1xLDvZOVIDDdUVX
bG3b7CL5w/BrwTyj49becPXeDuVlpxJ5Ow7e4gEb+arcP8raqcrxhpYMtmoWbcBQQebsR8B5qHbF
UuJfIW3h1fR4OW9hR381wWmaElNtqFSM1V6aYiBlFX5ww43m8FETDyl6wzTborwqo7UNYeOcXvds
wiS03ixQECEOZfrqOU6pZvKuWZ3GTk7qbQXKbli4OrNrkzNiWPtcq6YlaxJDCj+BXvLeBNJjKwwq
stA7iFyYfpb93OAB+mZfrEosZNlDe6fDUfys0qM5ZRUDYykUSCvZKewjK49tL0rJdbFdWPHcr7Jl
kF/nphXY8NzMPIll4/pFGpa8/8ltLoRC/zaaYH1soS8y351GXupCp9Lmke9JCG4N105FYvylXQ4I
1uqaSIV4MhyTzPxoswrV0+SB4pbfM31tAyovia2mvx/iHmByqoEyvX2LNUXLdujDvCgIgzvEYk3K
ISCgrG3OPxdDPnTyCLkwbdgL10bs2v/MHM43qw1j6a44GHVI3iFfdVaSMQGxVpZ5EHZa15ydTIeH
C5I38s/SenIacBu28bHF1dKwkuJF6GcLz14EVhW5k454CLbJ/L8MIycZfiKBt55m6SDl3ngoclby
yiVgTlsYwMq8TCBbYBC/7dltYERYS3DP1uVYIfKsn7z5J0lkmGgat1ZkmujSjiPmv+SIPwYODaJS
3D52T66UHNmoyvtMNRBXC7K1Wmw09/PW6CkWXjnEbFQlihKMHWlYTG29EabyyKDCwXFSctTVrZBq
tBIyvAl4XifOqnBwJMlhRoMWgYEcHH5soNhJzIszZIdaNzlUbJGXESOGTf96A/jOVO7EUjny/uN0
A/cMEeM/SAnUiMAledJhOPV1N78RQ5aeBGyE+XrKy+cTdJ0UY98EGvx+tIoW8fRqnrR4fW7fu2Xl
4a13y0uifeRo0+2r+7WkteozcJtNAPX18E68XoKqk48EDFN7DJSV2sIb8JHMEvgGOoKeXsKywjB/
cVRTqf0xXHPhIph2DZ86pKkNU8dTRul5EwAgXBy8iVKwcGX2EJFNGxeD03CZpwXwctWu1uOHjyME
sxgyDv6hqYZV1fXRS3/cKS2d7OPualv2xFRsxDMS/XoW3iEeAhwdfNjsrd+bGeTlI052HZK/918H
1tkFgv+m7kTcxgJJRc0JbrH5R7FhpyPSRhx7O2rh55sMdLODmW1uhN4Ib9lHhYKjEx5kloaL+FN6
N4RrAn1kpcVQt+vxdvL3NcokZIuhg/DBO+Lle/RE4riZvuHnqB2I2vbhRuemEKEK16NwEDAE9fWw
6BiYtMX0tMbpdzd1Jxcnu/Qg4PTZdjhuXkitBhy4lhd+GFtM7fhMa4YMTKCANrp7oajpij+nhHDs
liafnqnH2ZJvl5tKX3MEdvAw41dfbWvnFC5vfQ1Mx7wJNCljh12hJ5JFfMSQWG/OPHXXJkW4OtEA
PZAPo+9pbYrEzLH5feGTc2yHIaVbi3sFOC0jsqhKw3lNSoSKqfPRPgdLiUMd9ozfV0tyOmWsYZrX
AfSpAHM8514skw3eUL0tmYEnlXbzcFAcHSiF7MRYGSCcKu6nv19aR9Gl1AK7YZoOgEsC+1QGWPvS
wj9bgJHE+bLgnBzpwsNkzOdfaUro4uuRDR7vQ3wavk7g6haWAqrRs/3RYCBDMvEXzxjjIGsNm90V
xMidUk8DHvG9Qlfk3mbEO620rPE2Q7yINMxGgBwcHhLCfniyJhOOfqqRL+FfwP/4iRuIvI7FoWad
0VOdk3NxMSYaXmJxZU0D18yQyiFKF5QmsX4Ie5TPELX8b7EfynQ+sJJ+biscdY1j2JeNb1Y9sDi9
fagd+QWYRrM+MsAKce2JcqomN50wte5W/XWJK0f9rF8hWyzGG6d9Z4evOF1jag4m+eK4hFq2HEci
Ue+ribYCqvOkma1FHFXCxuqwGnsyQcID6+uxg0heWItjCmigjeYdQlRdW2y/XrFo4CZ/rkrGCzK/
so97ghnbUG4mbnimaqbhaabcWAk+oOLsLB61l3sLcCM9jwPpQu8ocGvnkSAawumyNEtibgs4pPMn
4/P5/QcdgkxIrlsa7pkHMVEbN+FgdYmPEqvjhWofA6VfrACP+xS8HFVDyuKCl6iTNCmnU2ep756A
zlrWUEiOVaNr7pVOIn1wnkQgVR/iPxxgBjkzcdg/Dx0gQx35qDKHmgdseNylJ0j9BpJsIfikpA3s
C7lPW/CigO9xzVovn8e+YPbVaMogCqlBrqZkNyHvdVmQoQQRX1QJgmeEKYCGzP5j31+cM/8bfv/v
GdbuRrpofZjAdCYpGgeyicfthtDxnkqzvndBkuTFmP3+2kiOp1PWldcop5wNuwqOQ1gR/Ns7tqgm
eomBRWgaaw479PCWGvQP8g+bHzJ34mkefC5HsCQKqaR0UOhZsNwqTjMDzbtjeSRRK1qUZGdOjLr4
nqbqvVIODFBO9v26Gri04NqcoIMcQPi+utD+gMw+ikND/t8RyF02RNsXIk/+x2VLhrGYSBrZ6VaB
UCQxk8JbMfs9Dwts7ntzmk8N9YKn/l2cfz5Q+PY/c3OUh0ASnFkldEH4Ob0p6MmT5+coRhgpIx39
O3TJXdG2GNdBkea5jHIKrzzhJzCSgMw0pGwiBFBv3AXNsccxUPYLXKgqxaenMKwjJXo2fft+SrCz
xDJGCxBJ4V53I6hAEJZx/Vv9X/pnGozbRrcn4U/oodydiON/O/AJKN0vcnh39F3A+J9iwaxvXTVx
Ui57Idv3KMjOvU+33JbAjQIIDi+zfwRaxedVci4vpiuV6+3Wl9ic4g922LAcI7PPYbhmn3/oqVJY
WCJ3/huv12ZrOSMjrpCo61ZsNHHDgGhNk0RMeaN8Z3aH3Cp6VgqKx2icsj7NWJh+5ODkCxVGtZS4
HqrTmVZJsu30wcFG97ZHaQYWEu4PF1tci/mf93keHySq9KQbx5ipYnAqDaaVKkZk9Qr/L1Kzl6li
e4LTHXAMnbNBh2Y8qCJjqW1KSg/5TeylxtE+vmUTlPpJCsp/ajJrJCE8mzI15I5iiTuRtK+cL1hn
0QbQ9587pq6J5RwjP7zgzue5GTUBvdf8jKw1hDVEpWMuciEAdBTG+2rAW+3BJbn9IQKx6NFcjdWl
QsZsMiue9qJtQWNexNH++T859N5+Li03Z6fk+7wuj1eC8ddxFmrKtIoDwRgIR9xj7OTsyWu/2c1Y
XHbhYpMdXJUatd5WXujF3tulZygV+MlwO72j7CKmpSEaoD4MIeoX34r5oLGl8k58d0JjSkrpRDeU
X+pRCL+YnOf1c+NLVleL1Y4HMOxiiF3ViiAyWdOjc0x/mjQmIRYqxRfafKqEPhZGQ5Ocj+wdXTcE
FVPrcaLcrAeY4VijwZD6Kt4JbzjQbES64TUFSe45c3dZsEgb5aICXngv7pf/vOYCQtr6JGSJkyqC
MI9cIcg4rbw7jVzGZ3Qs8N7FXOaZs+kVJHbsv+iI3LJnhJFgfxWNQAizSiLrCILJ9qC7ewCYIc4x
q8usmcH3JyOJxaar9SIJ56kM1K1gaLp1swPImuXEzfDMvLq4v1x14M879J8mRbNU+wOx/7yEazYc
kJbqy/LSD8mLvpTRzlWY27mNcpLd3kgeRN+cpIk13nGHrsPdRV8PK1HYzE5kbPW+KSrUgqtc8fm/
qP//6MascQNw6gGDqY8r2oTikwUYd1f/Y2EhjBKEFUe2EN3yolW/C+bXbcLdCj075cu0UoKSzu2i
lZ+7FNYNWmF0490fJgFaja5CGbrY3tfTbfvX9Tx8cSXscaqrEiUetnfmT2K1tZ5mPa/6Uhc4W/L1
pHxP7XEAqP8HMYQtdQkf6aglj+sr/THoei1ULrUUr5ZRT5XQwim0yMjiKLZ8j17hGnULkNPIzWfC
1TaKw9nQsX9V8oy8KZT5UBDGi+Cel8A3LPfkuaDROvH2GkkoQWtPGK5SmsNQkHVDg10hbjsMeTcT
KGjYMzZF7XnjXneqgQCwsIALayVxLv6kVO8J9eY1POHGuMAWaGQ6gdkZVQDp2Zi1UCfSLoUNRYfz
9RdQl6QDqEvFYbFCoRBpg28g1hDuAkJPR48QU2f1JM/tqPjlvPSDUJxAMAItu/XcpF+s/f66r8SZ
7A3+Xm+wSX0FvGsPiiWQCZucw76zpH4WvrSEs2+UUX9W9w8h6eTu1cdu3+boczcVN+0c4aBCHON0
RJsW7uHV6wKpxQCKD9pNPuOjGHNNAoi5E2rEkoRAynRKddk9eVX3KGlL7jzcRRh2qwafBKZO6VcV
lddrGw4unEKa+hPwfbY5YMsyyyYrjhWVt7TnXnFcP053r59R86paoyxrouirBRxxbluJwfDYRvcd
26aUNxwHgdB6MPy8HJr1llj3eIIKxQbgC2GwUGwuQroIS8CKZVCjMUgjkK7qxwNJCh88wXfrS9GW
VS6eXJOBX8psN7fKwngz9EvLIThEVRuIy/jSET1F+U2hOrXJkGQiSdkW3DOhl/HIb0eyOsf5Z4ki
nENgDRe3Uao3kPNym6vyX2HeR2rJpjaMH/tRXaE5np0zewONnqCcyOoOENB3+ZU4IyBCUKb5Qd6t
FRzOMWbrUOxaGUXG6603gLBzbqjQrzQimOz3+i2CWdOk/EsGjOZLG6r5ZCtZiF/XySlBO5LGlUFF
5hUx+TcCNKJGROlvDPaOXynpxe6tQ4O5+hHf9Sz3q2EhUkYM6J9V3Er0vEPZYc5TZd5TSairVuIR
CBtYUB6rPGUYIBhd8XQ1JbvwnYgIQjyC2v7vdlwv5qF7Ka4jtGjuBAll1wEI1gEXYQAm7mdPc9Xo
57a6nIpPakRh25RJqMz3VZMfoxBYgsYGAGxze3RAOKYZT2bjZpOF+Yy354aSmsGvTwbMBe74V9E1
0wmDdBnnB9TjpDdaIhTcZDYhYlrKUG0ZdEsB7ryvxZd/4zAo1mc8wFphEIAc6/pyjOCN13ME41Xf
E9j7F6khcRkA9tR8WfyJHtzSkie2SzEmvUozpJKZI/lgh5eY6ABHKo9g9BSVMR5lr3eZbE9YTKh+
nHbntJdO6f6CeXDFhutweD+W1xJ3Zae+dTmyc7b+PM0XekRAeBIhjM9ruCi4hg7Ka/Ke4ko4l6bS
X2uuI3GgHhy5yNge11dqnO2F6+EpquAyW8BLctnf0C07jkluno9xcgQLYHeW/DGmYqihBPaeqZ6N
SVNKff2xO3OZoylWoWDdUK7/DAH4uT2G+Efh0ABXAUk1XFowL5tdCo+r7VVyUkYtJpnEGl2j10PS
rUdiDOytauxkpgZIp9PNOZ5t+cpmKyya2YBBLQJDQ4vHUFuSMkU7uIElMH5D6jujfpCHYnhrCmGq
JuFwMbgowR1Tz6giqD4iLFxWp1ziFu42ISNq3wifa6hHDa+AczwwwV3QIUDUgsfxnwB+O12EK5V1
7SAxM3fvAHiHO9QGGZ8uHvbhEcyUfaZVQYB6VMAF5OAVANcpIv7rMICr59BVjP3uZIdJ3XzUaFqs
cnoogYFBFGjpL5CmxvIbfyeqG95JGgIxDMhRT4bOzYeqqojRWRrup0LfJavFByZzCeh0VTup/bNq
5q1hipQJNul1gzZFX2qxm39jWullolIBjagfxVucIzADlaK8SCEAlTB4oIJKAevp89kWSAr4sJfb
EfOMEgLzNp3hBLJ4+6bTsW23TY3ySBWcqOY5oOVQqJQln0gg6KqMTH3C6ArdPLSffgeZGJcYXUW6
quQNm3Qu7izP9gACNhP+dKpQyRMpJfrF32PRt8kJcpnxDmB6DzDv6QCXWfRa3QJZEqyomGQP1Wpr
bB2SHH4bCSbePkORyVwHgeo+RARV3A4+v+4Xy1UedU9IxKyvnsWZQgsP/CX64M6wQXh2mlj1y5V2
vJhJW6vL0P9gNJc/oJEmriTd05JCSumsvveis3p/WDRDKjSqWLG8scq609BL+h0/eY3aviK212wl
coXDNXx3xnLNrOKZzxTl33/yng5ekrR2P+ygD7WHad52z9RSuNHH7kq6RbdJuL47aKB2rT9r8prO
xFYZW+e3Fp1RJIwdgMERtix5esOCNpfEmWC/gg1INamb94/1UaUDe7XeL9UpT1/+OD3zfmr2U585
KZCfDPkpzCEKaIXGSN8U7if2pmistN3zxV6xaIMCvaLzjvShxSQ1QEUsbjEDsz92mMGxdO3llC0p
3TlFmjyn7J6zmFc8KfU0K30sOOihNHfA022f6s+TA9nbvIAN/LvYcNznTZ+nJxnG18P8zaorVVMl
Cfl4TJPZUIh/lQRVWZTgtTK8ifHUbVRWfksQhgncp8g5Wf6zpbCA4uORT219brHMpntIBKGpvUE/
nivPaeWGhD7en98Q3TOe5C/GNntNViKFDYO0Io6QWAvb/O/F4yKLUfLAMm2pBUO5G6AmyUUGt+/P
WGn+ocsdX/3QKmcB255bsO4qtOzTMeZ9MR7NNNvWNaPs5vb0LQPOXb3oraa/Yv8VDAvxq2cJ4W9T
7f2KAQYnLJcW1OBUbRKbW+0iLauLvn0u2wFW+KSDsYXXy7r34I7VfmOpOykCkCZqWNR+kpOrhN1x
wE9GoJllY1SPWOlRb5a5fUxPULMf6xxGhv/nVfpMyZcDIQmUqy24st6dsofYT/vdWTUT0C6lI7tO
aABBFi273JExAfTyHXeBi3XOwQN6p/HfdLP/rVT3vNN6hlinYA66/zPm8f9IGaE15bllZZNuoFcR
Mqcf5D/G/7oxjrR69SUMDOJDB+ZoEy9J5vDsku6hl+WjAyDePZFrf4DI6I7gv3m9AlgykTGY41h7
5GUUij5oucKxCb5eV+G8lB499UgIXuNhWKT25no+Z4DqYc3SOr2bl9kmqjFph+p6T6OSfwL4UOpn
+4Q3NDvpErMj2P80HwEKrFFKRsJ23z8xxC7L1acEhVuHc0/kKqGbwAkDEwNCUzaDQORCgZjQBaKO
gJMXKNyA+6p2qUawB7uWSzYFBiHPvO1TO8mgF8ZUvOcr5VfHC1FUKzPKMrgi/25Z0/SHlKX8yfST
SWMECBCmKeATSYRkg4g5K8m0T+fJjEfdQam8ksOVwAGrGnR5mAINsYtzgeLwqw5+scALeIy5bWpa
QyaNqhnowy9JViYe24HGwEi01upPH3o/lvdTIuODsr8NCjCUh96+4lCDeXSNvJH10sqzrjdEov9h
TCz8OuLDaCFp7lEPbhezyC4MeuPKsCE+seg1kFiHw5ntMth//ilC/3seb3OjTE6vpUs2xOYx9SgQ
ud3XEj8vgDWRKwhynuDQ4A5vEWz3qQg/ui/KF4v7bNgsKJhpLEidWKHWj92c857nRr7xTNpoFDk3
6YeqAeK7gPluYX0ksjwNd1lotBy42zAQFdIv6ZwreG82snCyq42wyG0eTjaRuExVMWfJH20n90/y
OjEMfa3JEVsouKdiP5lmgr5EQFc0Y2/0QFpYS5duQbUlTfc9e2zCN78v5RVKTnkaXN8fSuVGlVwo
kKQZdWbYmQwKzodw5T+9pvVBS2MHj6DEcXdJ2wrgAgjESM8BRnWu+/PU9ieWZtGOyFxOaNfAEPgO
PUJz13YrjDJOcAFvHHB3eEO6+Ww/5oOpXyc7JpN8L43jR8TonS4n/AgBBMYpFICK9XzLZSkGphqJ
+CvPwVWTUuC7LS/sv+7zRFIkieakeRShoDT78qxz7qtWaPa/vlu841DlBBhH0SYBP1mvaPRceY1L
7keTsZMqSlpH/ctfqUVkmY5UccfGiSB5X1evSJ41FXx225B4QClsJoT6qClyGpkRyeV7mU9F6QyZ
OIYtG1AEMs9pmQm9j9dYj9qxuWRPAtANrOjvhQ2n6YqEFZWZ8usO49gERDpPxMXsaXbBMbuiY4ux
UDdnT8uH/yTBWPxT4nWMCJ/uAj6DjiKpS4V4pmKYVMURtf9c9swueoXL9G5L1pG1q1CQ6uGRx+9f
DRAoBq4kP2gEf+BZSTpL5sxTBT++eQs+ti0lyryxgq2XMz7ZT5C/5U+SEmyEzOtOikuQf4iLEvU8
0cAqxLRp9Ja7dZZ3kDIexCmR0GUKzTiogS7E2HtjNU+d2le1uJu23ubBCpssh8+1vuhedWoOxBW0
/2z3Hf872mLnGRcvhtIyQH/BqKtqUvY0ZilA6CcKAFQtWNbkDQS/uoPwKkwRQFzuF1ZJeUKoTSmb
L+5eFwkPw0lmZwpD7BiMbAbSUtMVk4d77+R+FXW2C/TozheFlNnKmyO5SNzmV+PyINzMCUOvRvU8
5mqKhLf17pmEjepF4aJJz258vfzmS1s7p/lDicWTAlWoKPPyYDaGko6sbAYoXl9YlbRoB2OJ0oCs
khR5uLJ5kLKMQpx89jD0RnwiaAC3d7/lowM4FuUrA7h3vZ3mx4JRDots8NAUlwANQIhjv7fxFD7T
7QF0sTGp4nZKacIxHVBRzF7TzX7m+ggc+24oBgNoFAdkDvIKN58E06YJPTuo043h8LWLvrJDmCoa
0H5fXtH8IwQXec4G/IzFwL5CQ6Ax/6n/7NwfKRbysLwgk44vPQwx97QffNIH31dS8r1+kNmkaUs+
JMJMgQmb8/2PTjIYcPGO1EDyaUa+P+5RcO9Da99GjpmmvHdxBCPl3xDkVEsLIDf4ACfYl4gRx5rA
GnIaXSKGqBMCWMmP9r5EgBBo3E7LT0uOFkV6FxgRiV70h+OSLhI1/8zR5X7aluiVUhCkZD2q/nag
toXvv7D8vZRPmxO6qwOt+OBHNV9FPXbDwfYZynZvzru9Utvg+pRIZkX2eBqGjOERbPd0u5pylpos
sT8OPYB+G7kCkudsGZip/BjdWgsj3113q9bQeA6cNB+eZF/As1c1rg9Qh5eO6fLutH/z2Lo+a4mi
JvNU3mjxX+LAUxEZB+F7XXmmAcrvsk0q5W/wkrRm3JkAVZ8dbmCCDBYWa1EdCH2kWerDGJAIU2mL
BVxoOX+J+x9w+4sDVikk3OjdPTYZ5TsY7Qt2KrCGEODcFLrUv/uWwIGp8a95FOqU7vC2CQC/fBRq
51iLp3eJKSjitPHGcIjpSbYxISPiSTxXr3LYSweiY4CLLL4FXCKPRPE9a3psmtbEyZVfyUWOWClH
3lv4Ze45A50mzDRzFbt4MN0GQH4M2gxDK4v/WO/XzB4Q4GyMRuJy7yiZanROqdh7XC4BVee6IREh
C79OMUEox/gYLO5RFpE0bwxZVSGJnGWUMFcAeafzvd1mQ5cTSwJZhJsQAANP29/meh3cxQ62SOes
DP9yWgW2c8QdTNT22KL/IFPC2Y5mh54aA0d/TmN1mBoLESjE3tbFD/B6vqH1Sl4VtMoUSpSfjIs3
i0AszYtQf1DGoLQDdjgxpPSMIJJcMw2S2hgdeQYs7+JiE7OkdMgqFSGNMK/59VpF6eQWVVCsOzL6
OANR1I+oXgTJDBWJ72HQPdUvs8F7SAsP0K60BlXohgpsoQbEYByn6Gr4z+ILJfxqxIOOF1TAFmoa
0HF7GnhCSDnN8kjOVKgqV0tAb2+0+jkuC5Mm9f91BmBmg4RxO7abpZPIRLiB+0y5OmBSEgw8LSqT
LvQ4QbjLDR6GZ7OQH77XF5FeMqBOXoaPOO74P2zpeeEpq5bW8KJP4qpFEqKxu3Ck0xdPUU43kYce
f+ubI1FSF0zH9BqHgi0oWkwVW/Zha83PB/rvuIrXFM0COKK8YH8IAPtfk6xRT4eyy5s+zXiVlYlr
Vg4B1M29LN0L+Wd5yV1aV9CRNidXau5JDmJhe5lSXV5xYR/agOrtEZG+VJrqiHZLcKkS9bNu+u6T
f2agyfC1Gfl+RMVhaCsI18OUeaMwZGx84SUgC57CZbZqLVzCfsIQ1SplrS1iCxawCYoJ3XcJyMON
fQJERXlhGoCheQNpY3Hj3i60lnpLvxq4K8Ah4HizlELs0HkeSc7VCJtbtPhkPve3GACCtAhYXNdr
0rZ11UOmyZBqhn0gyI5za1rdmBni+tsuNOVlc2Ra9pHLAO601cIoKzmoJCZ6khDB1E7mbRhk9OGv
3kozRFW6PooAUrY2hO43zu47tpgf0Q5RbYK5AaPMTYeuAqoeb9qHsoaquAHPMPNjizRpFfdMuKiT
ZB6ki9BrTEboxewgnfjc2EHFj/kjUF8T2INzuXsVDXwpy0wrUFOxuYrRbZHPugTPt1Q+hDjPe4RP
vhRUKURMDTna/oanAaDgh4J8X517BeIwZjWVfQVikCnoosV+cpX4wQL3ProBx9UrBQJl676nr9Np
1sGg8nkhifyUSif4JgfJAkRfS4RoVfadDbsrDcEiUcLffN+3D2qMEEO9iwpU8NyuQ0kRr9aVtuuF
vHD6bJPcARfJyT1wK3D4A0ord0fhWHGMj15kiWjisTEFbSd0MTKmOUGGa3UlC1r1bIUvofaw6CHM
YoqisHnRFcqwkd3KIvjAT2lNZvvkKynT/W2fTHAT6+9qA3GPzNBSp8NHlfUS4nqOu5WOIcTkcGjs
ZGbVrAyS7IaBxqWm7/Ie/Ufs6eTyV2BFZcSt8lNu+TsZWkFZ5LvP8IRF44fk2xjieV1XGp7emIcB
2Y88Ylr3YMuqbOtc2sQEj3dCzpAoQW4JQeya0iFsbscOQwsqs/TrG8zqRZjwAfBz2qgEQ6n6LEaz
RbxLUAO6MBiL5KxsPcVtb5K798rqtKJDc9toAcaKxJbsxYfht0nOFEby7AY84LytZicm+s+Pqgfa
W4Yth20nnxjTXFayNmMYNk7W1sKuVqPsXdDoujFVVdsaq9np0GrW3EHh/XWs7tlVx7d+Ua7bQZfM
b4Fn+Q+798VWeeIZEX5FM1P6os3KvU11rJL4hXWtDz5r8qLccOTAS60iMuDQerhS9cvdysp0slIk
f0KrYign2ZtRHo+9/mMV1jeLsp9YMB4DcSalBtbD/QAHx1/vPlqHLTI6g0b5DxsMH/Ld7FF+L9Rs
tLwSLNCHiG+pI8PHWd7KAoezb/5m99tNJttir+UkypvC5Ms/fAPeU7KYeOlMVj921z/U+WEb8Gm6
DkI/DY3z3cLNV2IeXXCmmzZRPxNKefMh/0CfD7Oo4jtq2/0NpWuiBZcGFvLXXshEYl6JSuRstFip
8SeEFokUxUM7ff8KxBaywYkAPdkRE8cbXjk57IyscsxZxnpTCmbhRhfnn4cnrCVySL56SBlJmGB0
I056YXB1Nd5mX3CxDdUY9JXAS8sjSePa/rXMMJpZb1tfXOfMUO+Tdldi8m/hmftbv0IohMbfA59K
6pSo6jXs2LjSsM99UDGKnxBkpd448YkRetp2rHJ2f1vqqeEUTc063MLQjCpm/7iVVe7By4bkxi1k
aFcjIxNxbNXmY7Uq/T9mBChpTg+sKihKlLmwVQx8gn/EWK+cB3bSIMyM8j70YJKYGmGvkCmcI9Xg
t27pKy44KEQEJUk+/uLJfgpLWCnoX7/mweXfpFsE/ahIB8lB0IU9lgVawh9uX/eWSSgbQDERtTx4
44FOs+JWMFwkhzZwokmGaiyZN6/Zi081ngHg88v/Gg+ddyPqhvE6lCwte8F9yT8GDyGXKGSg/c7a
Nx6osAnbhaUGFmwH8ZbtFGiL2daBGrgsbZlF+ZQQRsW+N/txT6tj/vxkDZQwUiapE19EiKzYjzF9
/qCR9HzR0qWDNe4W6dx3Xjppu/TxB+qsCJz95wAGJ2xr3at1DnA00EC+LYdoji5E6Rcfh4S8p2yt
jAUkPDH7Wd/sQ39A/mY1QhXxkCI21B6dD0U86hm8y1p3DD8FbfwbjBUlq/E0jNx+yfIzpnQ3drIY
tCtQj4wN2pzfstrovkB+tF1icqn7gMUHvj8Kb3+QIPK8qg017+EwySVYzyjqZIJnvrXah61DOLjb
q4DZ801Jr9wblITQA8RGsOtpg/RVLR9azKtCWUxn2bea8zxn16JpvAuK4UruKTsCmG9AZpdtcx+s
6Jm6CcCfVuOSPOcavieE9w3/5QJxol1A6lFAbGUuRS3jJ5oDC6Vu7juMt3UV8efX64akXdKIWMeb
X6c6/0wKfPwICYzu6Qm/oIs2lKXvD97qD+EN+KRGkTUoMIGzGpZ+yPtDu8NAq4DUT8XFHbxaERVP
KgG4ZlL9dlCJDb7pk2/hGg1ZwdEdO20TeIO/0rhxDlIVHAV7E742oQKZO+OluAU8RSdeX0yuenjo
Hw69rPBdGcesJvY7MXMJbnKWfMGW7IMxTYrxGWdAKO00wCf6Pp+Jnss4WJEa5+TELErxsEUEyvad
moWHf0/XZGi6lGMlH9tH2wFMi3YEhkmp1W0L+mvRUMc794VMLr7kKdoiIIKzKYXaUml+erKaLt8Z
ap63O6A01Cn++lWQvVS5N5rvZB/Q74oTVxwwI4migvQYmZWaEOFp7T31ZgifMa0dTsYjY3IsCt7l
Xs7sJevjRvOw27ak/z/gHpEp/ORcPefbbPZNFly8YXB7zsDLYAjQGU1T/7jDbNa1xOKm1FzpaT11
tah/9eN35kdXACoiOQtP8YKUXVT/gDBopYxUF8FXKtw6AwWq/VnP9g0cIA/Gm4LG9sGfMm2t7J8w
+Lwr42Wx4UO++agVGIBS5s/ChOXp1T8WIn6iaC2ebkjOtV/4g4V+foFgfIokMOIYnEckNCW5WQyz
GFk2g66iSJBFIMiYjymGs+m+Xke6oZpcvrj/bnrM8PE2bfKoDO2yL0jW2BcjPoZo6WWfYjEIeJYj
vUHoab2CNm7qolA0HNy5dYqMebybSQu2r530hZTIObr2Bx5twS0jqVyJY7BByfdsygSzOy4Mmy6w
ewb0Fa8qg55wmlDBpAeRPFKYYENlZYzhQ8G5rk+pA2TCAvLlgHJo9idB0qlPurTJgUx0iSm/L6Lx
3fCmUnHKE1NcY2r9xdy4XFOQljfYSRXkukV2nAz1HyMh1xapDmxCJn8vCJAKo80IGJLkqFsmR48u
cpkzpPyceIWXkgi5GxG3UllYKhnCpQm0H2z7QYcvq9mDerNLylj6bIW674UEBc91PqXlX38G3aiw
SjplooFmFJj4N+o4O78ThG4mWdBjOvEjMC9Ruxi9TvAhGhRNcM3Fz4hnndCMAMf+GRgqMw2MZuux
bLXSAvZrF5MkEjkR93BZ5xLHMhL/UsEw9rq/AvYneseo6tlm8i44UPvCeMWvRu14qgz0WKDq1fgj
24qyuxw/LN2xbSeM5ReGORLPKADrOVGunJ4IF2Ta951LKzTnXQWwIZG1QrDwwxr1Albn4Ps9Uqa6
7MEzDXEvicjR7qY8/H7oqrKKj9oqX6au90ydJ3La4RSIJFPXgkByEAHORAqSwojg492/sJgVRzqQ
IiBVMTOiBaTQ6swH+iwmh5PjOVF1R3F7znZF17J2DHZralITTEeS2ThSF4afbyTAfpAvVbBqllK6
ChyOynn2s+K6+NTbsX/yv+gyDQRMM1jGeN99hEJLeKUm9IjhFoJo9unYmEwNPs3PJ88pXDvmKWQF
amFrHyME5VYwO+QNMYjwwZC24Uk04JAaOUbgzSXD1i2ASyFibIWY9+DJOxQvUq+BrSfPKzzRwmyX
yo+yoHAK5ekN0i+h9flV2jwCI7w34mYhtK+ylsBbA9W+iKtlDbopzbG45vB6s+4YNb5CeQ0aMLeV
2Jpgn/Jg9KdttzC/iis3Jj3+U8u9dcfMx6cBD1MtgpxK0/waALXkbTJVMjyEF2C9rFdWiPqqpTEV
6xxF+4sluG+Ewrtejc/9wK6Xtj918xutcbFBaeOf9SqwkWwLOP7M4OZuMARz1JaYuRXUwaImASxd
6rhTK1rMM38KD3v7Fk9KDhP/nWQaqudZfr3nxQNjxvGKIDArJW5TR1SCgEPh86PdXyJAfGZRASii
TT78HjjlWv1SOWXTyzPMenG/hZtjxGBDIpvh8GL/4/18K89CZNtZcXfeI9ZK041pxzF1NxAddgar
72ftj6yEOTCS0gNl5VCC/Wgk7uyYj4Q+fpMMj+D49RF/18HYpvCYJnlDjUCrmN1ET6VkPST4ErSQ
iKzE+M7HDrC+A34Cq6XmIjzdXO4ckgCtv7Ue9Zvd/WLZQCt3r7+cpV+q2EZ3GS0mQW5OZtEwKcXa
a2hs420k+amavkJzCRB1vyWW3twClWrGaEjkntPczJuiXW5cG+i9SWX7J41RsHn2KsYvu5NWjKg9
vX5gjEVCL7qyCAL9xp+m07kk+EYuWUvVg2BHyaExBTfo3xOFIeUXiHLAFbYeXvY/CqHn/H8TdWSu
RbYeVPUGEHsbeYrbWGcPhU1K7GTZLazC1SWe3bus1xQwy/uAPDlt8BfYVA1997q6lHq98PzJeNmV
mMnbGDeYA7nbl/EmZxsvbBXPVsryQ40d9rrFRwaF/jgqn8dJXm9IQ67ulXFvViBGiNGKEocXJQDb
83kozeHsMs4CF6S4vjY1RBb2jrP97LsMqv1Zmpl+EFlmwjbBSO2Ed6KMN9qVaGVw8osTZA0e2JKh
OXFUVohEX0U7NCIUSe02UzvDf/A6+9rfxub3zdVMeVxpXZUAFK8WCGZaIZyu6XQcYmb428be17rS
MGvXy8J1Cz26ViQ0H9xptxbR8XUFkAESHSf7/XYZ/hqkTQ8OeEhdDPZiCFZ/nxpWnPavRjyNOP2n
S9k1uw/VN4zm7gUOSdbhOOpQTmun9yASo0xB/HBNmDBawum2Ux9tpF/ie1TqNkv8rj0dKNh4zNZX
pQkY6Np2YKKXHrcZaQkyMDGWKKRBUdxY/FWhTEJn8SEwKthyLy7Jdhkd532DShkKbx4VvsqRuB97
HJ+DwftqC0ku2U5RLWUBrf4mCAINda8pHo6ILwtodXf75nRGdNYvl/oK1YJmW0z1Kdci+Tx9lFmm
nV9oEbUX7Rv6TAAuFBVFcHA8Lr8nqniwIqhjYGSqpXo9BrPMJJxFFOaqiKKI8/8GzdCF/p/0j1X9
ZTRDxyp5KcosQdtc1PZDvI0r0hNEQds6CoraSPHFvQdzLji0Hpey4lxVH0z3/NzxOljpP0JDSLhZ
z/wihuoup9l4yYppPl6yyIhxpGWIxO2w/EQj7mTdTP1pNkmRheLucu5vB6dxL3giR0HSXkMbDq4f
lT4vtl72MfPuLd/6V+IUtQ38NjYEdGja6/hSqEL77feplZQwiM4FjbWiFKIKEdGhqzRPKt0VqoJD
amfEwrLHOQtlhqNRnaTLwr+5s7MbCfi7xZWHfA4TT7xWpYY9x/vluPbcOt6gWyeOItSGsCXji7zV
GufIJsNxubsn1GYBpc8Jim881huKlieBXYQBWnml8w9j2PTRrE/JeD0VUPZqVfIJr6VCIo0cH8ZU
8uIavoi+fs3WmLe8UYnRL7cjF44jDE66JwWisK5HLVDIAiEoHEpHyTL1JUwww0nzkDxdQeOYBY63
T4HyFSVBrinVZxcGPvVbVW4CBeEjKZDrNAsc+Ym1uJCNdIOWTq2g/QfUq71PRYtvNI1/gvTo581g
o3345M40wIHg852j2ru/HcG1bPyKyOAfQ8vWnEI2HPs6R9PAqAMzzReGEt9+SIY5vYg/7gwWHQ3u
pBda6oFiAXyBuY6hrlAR1UnO06JBu73beotVSVUvRnxQTGWLZF03CsGepx5Wksukjh4EKzQppA1E
QZgYai4ykskHESTzS4WrWhe8rTay/Ofe23opwpt4OYMaw9Yi9ej02vPDdoCS/XQLljENPzEjgaX/
OYo6oNKinhG/opVqlFe4CMGTqj8yxy25NA/wKIzbwd8k55VDdKprj/y5/OhzmFsi3Ra0x6oWkX7n
r+K/ZHG+T72tHnbfL0hcxwnnWA7e9E4xqLRqFbgXPCDssoAcGaiMI+K64hYYP8ZbpyUKoQO3VwrC
gTlH06cr5r1S6ciF4xz775IH/LqY+bQdYEDjfggaN6+un/DrK4EpHc5ckjRnpG1E1jKhsPsn5WEA
gUks3GBEjpY+8rpfuX54qs3P+kP6Ev30C6wCTsahJv02SI6cKhXXy9wfdGRMJByTywRHDSfvIh9c
1VTpivSKpI4S8E/QfGA9+JJBTSlGS+xozWzoZm2J30kBBsSqjkor2Abt3AxGSXg1RJRHMWBmL1jN
3kYb7i+YG93+2sMpnf8W5KgWWhBEIeKQZcwLXwCg4XGdeyS0VXvY3uPo4+hdT7NQ8CNbGkq5eN+n
gvqpxdO+krXTGlQ/6ieWawFuowXqSVmDEe5wpQbUc+41o+lq2kDxV5hs0RYIFwV0CY8+BanW7sRM
V7Jku0ocHgO1akqEdYU80PVbFCFmrzl5ogYZoZbTqaTMh9fG5M6w6iwESUIGltkA6zz3J0fDH49n
MiqXCgIQb7oudxgJhuzebvFpWxUmLwJ8WwOxEjt2OKV7z0co/nnPMk3c/4gQQnfdoezhEadQw/ZX
CFP/7BQ84dKfNYbGF6mEhANLprIM3M7qSnNUvPauhJcqPbvK1UnjenoKpnVszY/wYjNSaiMx2GWz
YMJjDFGJI/aAzVQl0BuRxbUObWnAix91DcyVvrA3jmgL8iGCEZls0yNhJBkyvpkAGbxVYkxLIaeI
ZAVe1pqWPnVhMTGhVk8QFTsePCN1Yo/SxshYcUjkDNdyvhcqytyPcPgQljC/6Ovht1Yu9/epbpk8
EDgP2xPnNzwtn2fG4cFadYOs5+tp/4GxGZGkT+g5N1R1CCMHHaBDyglmdAZKsXpfBlUAMyJXzddL
illzj1pkYDBclsNbGjMAA8YLyEoQUJCPoWFkzlxTni/HSQXRnVKMgyCTWiTlcBhS7y4+MnST4WoT
tpLzxZ47TNOIvrSbQ/Aqp6piksSEvf86xGDJCsXfxvFRimuUoOaCXa4vAcp6EGrhpovJSHOhJZrf
0pUPxxqt6LDnHAtCg6DGvBYWVNs04OVBbUDOR2y0OH4nznFAFndL12lkIoF+YmuseDJ5c8O7W+tS
noCzLNm8W3wZuFgh86F4RWxoKP9k8Mu4TBkiRd8YAQxZTjbFs2jJAGkEkmDBayN2c8vPFeKClfxE
PXBBN3ck1ssGMu3Z49WTh7locVPda+mLuDeuU9O9w85hCrX/vInC5QnZ3R36hOLtNu3Al8YUivi6
tY85WxqqBckPhnDtFUQNDFfQEANaO7YLJKVE16qPXhlTwNgnFQXIdAzKs2ZeH0GHWtjACCv+dqkd
r1Z6eaGt/NiEG2nTCDmu96aQD1iDcAopDDPg88czlC8OgN35VxfyvFpOXxg9Ez0qki6jBHEX6bXx
eF+mpJHrczhyWm+Mbdk9fpXFzHmHdlb8pYqzP15h2q9FbvIe5zCL1BnGbzrX6Sy5yLmedUms58fj
Ul4WPJ8HfNATnYaVf/pw1SbPP6ehtTdPulScZg9qrBaGriF0W0F2UhuoS6SdPtLNLDcCqELc5QVN
PMbDmP8pSMqBJxM9spFLOlMsqpnKEnGkdskhNr5notIq15Q4Qoy1IzicJoQZObvWvnYoPPT8MlGv
c3OH7bF7zPXzOXdiUNNAvuFuXeT7Vk6TIQGq1fyZuufAlQ3r9Eaj1KhgcZSs067bojexlAmyisuY
cXL9G+6CZWi//fMwcCzinlMSFpsFCT/mDHF34vLFqolk+FBR7vJ320OrxcCKs1w0K70x8JBBP49r
6XYlPb7lTfHxCvkkWHP8OcoGazHZ+eRsj08dgwjyYJbQzWAJG++EmG3F8MXO+eOrF8G8yolMNuhR
BET3iaHR4+Bz65Y+kybgnyFPHMhYBI2xW+KAPaTHSA66VOaBoeJgCixq/D0gKDlKydgPrPB7B9cS
JW/GhM5IAf0gYvMD6DjBx7JMeHS865kL3EYy/YMD1vaA6u6H0xSi5O90Kv8lrcXgbU7e5vSGBspd
6LGfUCgFVJKBLHmoZlZ74TRy9uuj7rOHbTQ3dvZ1pqMMmrcj0lVYdTVipFdeCJWw6heCTcqBWq1b
32FyLHaT99DohcExgUdpHc2/O837CTZ6V3WMoorb71ugQSPM4yfcZLTM6uVtcQFvtHFwn2ES00iJ
kayXqO6y3agV5FfcVpky6YKqhMWVcf9m5n/3KqmnhNyJZVLGqIC2jnLYY30lCUyKGk4N5Mgu6/lt
oAWo1z4OCqsT7KXn4QlZ0wEFk0NnNioptJ2J/9bFq9nGHSSAj6HV9eOOjsEj2V+UkLBvtdjeImqt
a+WJ9pGIQI3RIfELz3JLZtt/yXRka4rZ2+Vk/ELQG/aG5BhqkICIjMPr1idMBhBBRIar2N9B+c+R
YWcvxTCwu/KJz1h01GM+NUq8U7s0tqGlWu67adV3aUnXq1u3OZdWkAnMPxuWDOkIObGA+mnrFK0u
IyDCcvUCiM4CtynhvCyfOmX3wYB8r3SFtuILTv3KPrnArV5ZWRrjMzx6xXJO2o3p/9/H/rFxxftj
EBlMzc3PLo6Pz8lLX4i2KjB8IdPvCGgJlG+Eyn7yk0DsJ2GlQEDf87zwhL9+Y+MXCV92AKmjaTBw
Q27wfenxwXXZc08odpR9i5GM8Xyj+7G0F4XUiqgECfqYKV7IuaImAN7LktjVWOitdRg7EovjTuff
yXbOWqSXl/Ud3IPnyOzu5gyhjEmq7bHmLsrUkvELZVvdDCxkxhn2uPEjfsb4ZzL5W3/5lQIaU6KM
aOwv+yyyRn6VdEaKG9slkRDakEgIBhWagUWtMEOo1gWeoveNDne0Jr6kC/A8XioXCekxqEQ3EzUC
kQv0+/ybfqn2pueDqoPUDg+aNil8Au77D8UC5yuTX9MTnhR+oLgmhzbVLLToVZ2cRwHVqSOlMNX/
v+PJrKTZVF4qUdqqAdpnhZ5J05x+XGMekl3tztEFWRJBxVc6MxjD0bg6j9jvr8+jL3GBzVTwpUoX
mCCewkW6WK+oEPKA3cvCiOa6wSzCOL7NruoKwfLbVxpR1mTLy/Vvd1gA1MBNJW5QVSYDHAgBW1dt
jj02w2vZRf2S8zuCxPnrdP9gs8mmQL2VWubutimkQoYXN3EdO3E09bMNK2tAdcgfqWPcbiM90Mmj
zwSNLTOm57BCBcWsciIi4RmDRx7tCYFUkxHnIyfRNKG4s3+mdTJt+bTzzK4Z+mk0rm2IRbqEHXOI
G8vdFNsFuEVxGSAS7KRTnPTJQ/ZMs/OZWNdOFNzV6T0//BXT98ig7HXz/26kabdrj895WmJY2wjn
/XJp+R+CJ4PioAusEF6bvOCiunsGFR8nxi1BOADd7AQTRcPU1if3ggdLWF3CRmNJprqpRwIHsJ1f
DO8xW7mPS5s007D44apsiyP06BG0MnoO6Hb07R88j/ttMLNIcrybuwmB1YHFYyrQMq4d6GCn2Oie
JoADDnc+m8xCfKTJLUzpIeibzKm6uBg4RJnlRdUItxnOKiL6fA+P9guYvujtzBiqdHeVZz4Q9RSx
U7pPdFrji3vhkQ66aeh7TeGDR2tLtyVw6VhwB5bQh3wiqFf97cdwGrpDUYpXHcTa0H2ZQanZVsBB
ogJesBu4o8t7V4yUAFUJA7OCqRimgkGRuoif3S3FLqEqV75vogN2gDJ17hhIWumMjBsSVxI3600E
ZPdYyYaVt0jO7ezHCqUgsLyeY1bp2i4c1WAMNwIyWm1SgSZTx9ZGhlC6BGOgMGOb9kT6H1GJGLyd
zZaZxH6O9GutEbHfALu1KXJ66pdXtnwa1PrG2gr7O3N6vNExASZLNq4A4a0B2GjCHVlFz8PpjV1l
0h75/naJaKcwSyBoJZlD2FlaA61FmbLri8Q6v7IjWPNHf+/PlY74Fb478XRw/CiNNlz0WMf3sgIW
TZ8hW3a08AMipNBgRUt7lGN99mn3N26u5E3mnBB9hrBOOEgyjwWpAE4/ooALkJBM8507VIZM3hfe
uMQCQAf6Dn+FJ4mWLCb2CM396vJGXI4N0zmot+WykJ7o9Gveud0EHeVs3rxqqOUxB53XRJPh+uKn
yMHsSPucuHQIWZ0rX7+L9lFEL6dQUSEo7RHsLiUFR1+T6QhIRfWli6CYOTUz+VL/HI1YE7qPknw8
Ic9NLQumJRQVkg+XyhJ1j3nHc2cRbyUJGwcqt70sjVKw+kgvq9Cyw96F2waNYMKg8VKO2nAD0TJU
7qsmwZuUTIPEYCHHWl2ORK6kk41Sr/tv3WotWopuzae8z7cadmnNpI63SKP6EId7PRgbo0XlLGFu
kAV05pnmMkyadZxIQiV9S9e6bm5FgfTrdPQKkbE+X9pql/JypYvnPAX+10AW/HfmNSRJsDrhNBII
val0Q3rxDv9NpbglookMn3LSx5rpzhgzANQZZBmVnH3AIPe+Pk85VnLbWpI2aI221JW23YDSGEjV
89uqnNXYKDJ9ALHyGC+gVKK5bOWMySU4nOULEL0SO6IftMCdqSQpIJXCP/pyuBZIgEmNmcQ2AR2B
yJCikjKOyiFnzxSs6Lrn7nvQy1zvQ4z918KcG55IcZ/reZOQ0wTzG1USX/ABxTEkIkSsUutvhYfu
BMnnorVOS4r9O6RQ7TAsrgaatipxZFVxA/VJ5ZcitQg/J/e9qSCbPJzYpDe0RvsGBwTXIntROxW4
UC+Ko6J/heQvjEyEu0PrnVZZfB99fwqWWfG8b7IySDgNV8znMCcjVlHR9AavcVQLPWPcWTg4XRFe
6P67Icy7/bjXRezVTbsTC6lsoC4in4IfPd3nxwZ4PZoKUs8tmgiJwoifWJAkmrPGt3SEnJEbymFa
QW7tYoQSA050TqATc+gInYiKACNNDoyS5eFdDYz8DOBXLoGl4bLFno51+5SWX2xLaUrFv0b6EmGJ
/EKCIQe2FpjjX6bkjyGFq6gMDrqbBlUgg/pBst1jLoZW9u+7jLwg5De68LJCDnDAg/wxvrju6IUf
gWJl1f6bJ6SCnoZ2Bs/TUUKNTFTS0Gbr7T6zJshu9ZuRP+tozMn8o/0HKKXjpVGmjwx7ZlXdsFKJ
Xq+hgaZjE/XsemIEyQaPXU4W7qCSHJbUS/qWflCduBA9732SOC78+vu6enmaBADzK0ZBDik2VuKy
NWJtH+DBVuEzN6sArqp0f7eGQj2rtZ5KJbLSvnmaEDnmSQJJdfXmlU3oUXXkOcT579p6p0sVIFkt
vKxtygsJNdpI4YxsVFVjwzxfxeZrUttMPVnuQTn4t9vDlle+821HWKhLpeA1btvlc41kyPyVqizv
1VMozfKV3j8rLXTW8wjfOGiX4LcpmNsL5r+yz5VOUsXX7rQnkwzCtFKEyZVUtEw6FoaW1TqKVO+C
wmUH1u6hvv1InS/qKooyP6bdvje3WKoPPNa49cKDj1I5EoDGO/IEK6zt5ohaXi8PrG+ObykI9n2W
/0ViVWdzfClpH9x7hJeGilcJHMIoXCCaSPMeC7TBBhnpyahU457pdy3mU9MBlzhkA+qAGQ7CZIdi
/+1h3Qkd1XPOqpaYKvLA4UlVHbMviqoo84OqW8bMpKWuFjP7QBrMKY6aIPp5Ei8k5qx704qLDieq
MUmUI6HIbJOBn0epWdzinvdHHSoQTHNy9U59iEK3BVH2owiTHYYf5yMCc8CIM2wUrP7jLBPuYRq1
rYXwXyKZgwMpmhcpAZXOLCHF6ijpXYHRJsFzgG68tFIF64n7wNh327xWDQiHelkSc8FZ3YDmrTM6
VByUwwd8TkXgpwm2t+30+5Ue8j0RdrbR0NPe0JvUc6hQ3W7BCMoWlVmfJpv+v+LaY7p3hTKRgBNP
Hgp3PFPEMZbE7+CFsdWwJsgHcsBN4utS/v0OMdX+wWoMa+XOnCOcZHi0sxGqBMgFyU8VtMM4EGg1
mKyNXjxgg5OFj85hOeOGsvSeV0LzFMsP/wWwmybjliXD9Xmb8lWrcYDUvuWRqOPsrUnQ1Pw0+O+6
HqT3WML0kRhGD6L8fdETKaGM4WNogG8x9QoXdd5UFT3NEbM3zuZzhVpHwamAyoLmJrW4yVootDan
eJZZgm5bEzogqais7d31/etNFntBaMa6enqDHuZnJBpfhJIAA16BX87+b27izM7vKC8UDdmM3KIz
B/+8U02ShAO4CzPE6BxdLHR9ykJNqlkobGT3CnVqayQkktZmYSIMSruq2uYrVbtyyFWYXr78j9C/
ArcSw4tuEVzUvlvckkQ7KoLi3GIbuu/yvVZQKwZce7tRUZGy+sY2DegoQFo48xuVRD19Hbh2089u
5L1RavWibRr/HNpzXN6IgWUxuVIsWVrq7rzFtfs4WVxGsmwjGbYe1YkzvOTITwcxA9tl8MtpIiAa
BW4ZVcwMPdGAtTYdZAN7XVgejiaqztOmtVEymDV858U/mfDTNWw+LDAydgOcw8eh7T6nlpGOkfqn
lG6bPHAKct1RiJoTcWACqZNLJ1ZD3sbKYC6ZxsgquxtAoEQhb0YsrssHYfFT1y7rB8rharkhOpzG
/GICmpCCHwB23eRRctVMg9FW0N3jBazL9451AN1zXCAi3S3AR9MZfta7d3wJUVhKBT6qebyX4YKi
HlBzzD69Rjbkecf6Rzo1x854CZjL9GnMAhwrIB6CfPItTFK3W00xBEf24c37l9YOxM4vJxcKBJHi
zerGH5fpF7NDjNfhmP3ux0wjQwF74+ojIMu6HHpPzeS8RvNmyfsJT8hsNgZZ6D2TI2wj1sb1oL7z
QAvHJDcGRxK9E1qeUldanORBZWvF6WBwlL/W8PcxdPoEeDzr8/ybgD0tUKW+cv96Nx1HnVjMLCVU
hPMtruTbSPTrw9vwYA+WbH/COIDVrMyYX6mcSj4LB0DzwDj312MdxhS6CGfSJ2RI3ydKG5qInNHJ
vZa+pOG8RZ6hAnYYcnJAXA+kTYBqTLRbgYv3RODTqlbY9VatKNiBdtyJi3AmXik3Rw6iJDhUZEjC
+ROdrrxCw8OQtgYhbDhAPVOEVxyvU+mibFzxEB/+ohhyUDXbE396GPfUrIc2il8+d/c/Qa38Pd52
xBoLW6kEHTi6U64t7HaczVXdkZoB9ply73OT4LeMp9XXjnICewbC7qmZafQpKG5dPmjBbdctrcBP
j9kpgrLyZTkulTYFl7DeFDuukmZyCo8W8CBg5EQ/mXiu6+iEy1Y7AdJg/RJvHFShXOQjsUaoyWw7
hic0zHAOq2blUBhr5xAIV3MVpdFNPVdMZJMvoyX8Ne72dUeRK8UT4WRI8zuKczMZn1N3Dg6ZaGTv
8BNZ2pacNearQ5Lnb+Cb36wvx2ejH/f+IUcSI8X8ITT7QxXciSbP19g4vx85v2BrdEmaHeljdoIH
YpD8klK0XLn00W8MekiEwTILRLpFS9kOYnoQ4fKrLVeUo2TAPZiEy5x6TjVWNAniYDybqecrd5++
4HzBGXPLX1uHBm+sK4ZfTkMl3vzWvY0ux5juy3YYdbaO4znxshlYyMFi9hVo64FEt3p1ZzI7csdK
pPSoqzWsZBDRSieeehU7Pj6Q30l543y50aDuyYV+cBQLMIrNVro6j0zT1nxkCV9QX08ONjFpFCQX
esblEReC4RUzN3dVL8r3itzH7XXlGeHWleBtCCo2awKnAqro6VcYo7rXhEkc/K4qGIzO6S2iavUN
1pj4afC9kvaaGq/yCxPgdz03gnS4+3zkHTmnsEut4upbZx7ZxLWZpry71yryHYWXUE9Mn0oCWCTZ
k19TC2Mc4uDKxp4/TAWnSHP6U425Skht1MN8mRXzqdlaz+vv9L5vduIOwSQ3jBvnSJUxtWBUyg/f
nzBfKKyDdUsZWkGFjIAz42hahc7KGK4/LssXHxwA9SCBYZjnlUGjaR0zzBx0X+KZD2o5qIGEZPIW
8lB93lnBJ59pfPkkF4QiEuU03Wn0bMaKmOIzVzNr/IGKF2+Xz7Qyc71LStcssER7HemdxwOcARwG
OO1crgXIUeXPwI/Sq7cIqny8BNG06mTeb8QmNjRGXBjBFEbEZh5WDd82DVw+90DZb4Js2XcQWl+a
HwQ382l3dESaJOHYYFbTYON1ZEdHylwjWe8xo3wiZZzm4IhgRL0usKCjVLCzzXYK2FAeGFm29Jc9
mJOxY0sWidhjHv7xQLY4v5+KOEbN/QOVN0Gq9+mVKX2BMCFVTStwN+4qmsxALoaRRRK63jeI6jgI
H6TALB3srqx1dA+NbfOz0nGMMpcrn8Dh/ibnxc9kgkpdX1Uhx4EvDZKGRvZL2FsrzkesTA/Tf4xr
kDStjXYtJKHoVnI+78/SmdygLJlhgP0RdiHyopZCKa3Fykyr4Au1f2i3VtLqolIo0xleCA5JPwgh
4RDbDJ83TT/OY9KlxTngqTjSY/P5vi15fr79rRQho+0NbpA22R0/EPlOYB/wQaR5rSxPDC10h/B1
JzrS7oURWXlqgTWjY2AnPwUjptuEz/GXhG+dz+vVI13iCIJyekYi/5hA7afwNyUweSQeN+CONLB+
QwAIMes0GDoK7/M7ggSvnMoe3GcIOGD3mP8EqOcFQTCtF7U4mnyA9/VbDsuBKBxs0gdlKkeS5KTs
gsNrDuCbk/7QqPiOJCEMl0SPDrga1jREserTuRExHWZHM62Cx+1E2IQpOn7wN8cvah2euwWg2mQO
3TBnTXkKQA66v0WXb+mFzeIlznXeOtgCpvhzPwfSoo16Ny9krdcpsinttHFEVPGgpp65okCmsBbq
b9fqQ+Ya2ZuJ7uMxlJT5DXDT+vO8AEkOui1+v/upBSzLSREwNLoJOc6PsJHrNPQGOXW3SWxIMIlZ
2NlSo4G/tbgVE+T55pJlIO+FwSvA9LQIsDlUXdkhyA5uha9Mfh8YL8/lIgb9ZKeL2uDyE1I0ILvo
eCBB1nm+wsXv5MezzPhrGiwX7dRGNQDR58FI7+47ZRwhK7Czpt//cfbwUaopPHBR7KPcizQ7i0HE
UROsrD4uEi4U1oSRRFH3q0vZmSizsmvRxADeZVcdhUl+0Rjy1gZRmpICquNhJujKfnlBvDb0k2WA
BJFjlPcQRFd0fKLoqHUzq08mGqN9U6mUWVYGIg8EoAeMOz0kbFAV4ABmTzuK8MBeLCzNu9KezAEc
iytpAbfyQ/5anAryT2otbyvAauemSOpiNc2ScuDdDTQA6BFLU6AxPSfoowE9DjyprrGX/Wnj2cUZ
wFN5xVgX3O+7UL48s+ky7GkZ16r2Wo0F8yiRVYbErQ9IIpfvB+QbHzylqwN63/n2ShU9nmq5w+2C
NAOriYfU1aEPu5b7hb+V+AWAG4sXZSz0zAndVqgfagWUtf5p92j/gwKRIR6bRs3PyDhfHRAEigGK
/qr/F9+PgIxQzA9KgzESeHLNtMo6z4bWFWEq6DGR0jqzOg4oPiT5B+QQQGUd//MrQEE+0RpujrjN
BdXM4zlv+ipel4x1lEDYpBTlQ0HuizhVe1rtVgB9lEi9HHWIUXYyOApFpdZHU6nnTQmUv+ErInTN
8sTodmaj6sFcfcZ6IMuukVLhFd5Oh5yVBq3eM4gckzHZYY3yL/8t9CsheL66WLEh4rPZRW3g8B9+
QnCO6zBD6AOhBrHdRYfZi+BC43ARI2Jn/RhphMOR0nRuRtlEUvzq7YksFrmJ3dm1n8eA6AgCT4lI
O3/n0xUdp8DXweXOow1uQRhpqC98w+qoR+6NM6bmInLlmxSEDibtvUdjtnvxEZIYGJ2bzvJPlRtR
mXuLu5dT5sLTLtH/F8oGiGBQ3SO36+mKBYtuTW6onfXqhCy/F7dRDMc9BFttoHF5XfibSB+8KWg8
xqj0UHy66+C8F37hoI9aQKWosyp0HUTXFLd4tbvzaXictcC03aHMS1vL82zksu4VSGNXGm2c0YE9
c7f5zBt4mAX0avmkQzb2fbjJLk5tZVkZO8LIJPBgVBWJcvNryMI/azxkjNfnyEJz71uOX24W1kV5
q8f+m2fkqadMvFjGrKumkK3i3EVAqA9r13+yAJJvge0+sh/KHjsynNyNb2l0AS6vwfXUI0yk3ZMG
jvRJ6lctPfURZ013p2AkFP0dPKp55Gacz8aPmeMl/CGbQlgW4u85Q0kG+OiT8M+c9uZRDb0i0mhg
NELkBHZ2oIV7+uPiZcNlzjWhvZtd7UvB2PDvSjgxv8+365O5enaG0LdRk2O3Cl0LaxBAMfDpaNbG
NT0HKyvIWoKbGjCVhJqQPWNcfrwiVxh0pQWPp4BX/vNSqTQuvkN/84S+08bVplPZAPhvJDnsjkLO
6AmBNh78AFzMhi74pwgMFXcETl2C9RpBlvdlrqWarcRaNM6SLIFLxATOBWaoObMSp8MFG1yMYrny
kxGw7XuDVrxpwD5FHYUmUIwWqEsYmDmYXU5O6O6AavVGm9x0qfADY9SLeo4yErxJpBWsIeN14JvJ
8bWzLiG2pw+RnK1m7Hr9TJxzJHaWWTgZ+0JETWQPCQxZCO5NKdYRpU+kYVqNTQrwP6jdCHcfx2Cx
5IEA3oSLa+tikDDcGoxGtj2pIwDQz8muJZFOuF/z4LPXQ1PWNlafm0jUS3GxCvYnIGmtMKYcDkHM
ozwcxsX7aLIbiEUYcW/ioC5t4/xPWjl88H4xTSor6cOKCUxafHeJLVhAEkJoJEfk0/z1l1larGPz
LslkNhLLlJgeo/JA6E5ibSlCC7kofRLV1VbqwKIVy8bGsmrz2RW8ezsNdKzvMvX09HD2jCi+ITBo
yBrz0CRD8vgVBsTBw2rQjGfibaUARbd/LYOjsIsILtJQQeVn1xtrq0esQJXUv07qIVhMCewZc8dw
dvkm5F7H24ga8BrXSo4R6BRv5dBQDFgps+dFulZrrCR5hkFcFAPvfwXlGZ2pwbL/RoW5GwFh1Iqz
O3svQeiXVMZ7dvXFS52lDJBq/UFyAzAgnpTpGT1KwuOAEFQ0M06636wKyCQjQDPA5auqLdmE/87H
gQrafbYdEuDhB/a8v6EGH4CFLZWhB4DIbjcXuvtOD8pgUUQna7F/Fg5k595FuVHffjdkMtJXWbsZ
YkwXHmGyyfSjgOcZtCnvGZ5EnLYN8r5JpiY7EHF2Nqa5Z4ZEJCCL64h0Ei8NnSvgtUIGR34fKdjP
irA0OsCpFjG40yhNGWcJA2gc+JxfUxdSA6GFh3vwz/E1Knf/jc4541NCAmItrK02irRctbcAL7pd
ZpJHt3I90fRv4KSlB0gWZh61yG1oVHKSFkhl7oi0AJX31ayVcY5PbnkGEO6PJgwMlW6nGXEJDcJx
n9S36X252Wmdv7HcJAtW/vIv5JzR2pPi8+XktIrDf3JFbP547NtcH5070d/sWDNlW/No5hZzEHH7
7I/B9x4c7V+z9pMedAAag94uvSsDJZIqCkmu+Dq1cXfJz3kIrT46mtUR8gAjILgLxFJuix11H8dm
HZRVpAt+s0kH5JlEq2sLNUerIwZ594o1nlmdsxWPro2C2EgmoIjadnfU1b47cVLDbgUpGZ7eKU8b
/Ow7Q9ISVFkGYKXfNnkwWjCqem9ZfmH5Sh8QtnEc8qesvyDInCU1Sj+YePgZPwtOX5aoDYb1y9ka
BnPFvEn5NgpkV/iZeBdjvs7nG+DOF6CqEfczlIOrxfMeIzZUZby2Hlox4mx8Sq2si8UPlBQ1oYxu
VlSXmSxtypVFalIVZL0Vtk7cfjNUD/UierUf+JK4JqPJd5Ha9B/xE8emvCCbh1i1GjtOJvRSGPNw
z7Z+oXrwWCwu7va9IkCv6QUa9tCS8QkrSjMqR1W4BQImomIrslwO8qURETvsz9LSe6Mj4SH630qI
HgzWswC3k+JHIflDX/7vGMsBiAXE1elAnzrGJEFgif1WPoHVklYjaM3FSLuz3SHPH4mZmlYF2phV
YiKW6uyi2iS0ow9hsRXDfw/PAPGGtHWZqjOjM6j5P6Vk854TrWkJWcjcpPlesFcyflZZZnfAD1zZ
dAAyvNi7Zgbr19y6EsLTDaPDiWVzPFRFsnBMmZz6mUvHQJ1Mq4qVmj6GU46vlWXKm17lCSkw9s+U
YvvX/vyhHBde9eOXi0U0Z185bV1htXx1rY8UtNoB+55tx1ztwUKaTkGH0j8YOeLhv3cM9Ir+I9LU
nydCplKoWNVQk4stL7rT3Q1QsYnqGBl7RY+9bgRQwX+V6Itw9IXUACPm7XFbnNzWOGlNNgpOB997
2DFi1wWjVrC78+Z0OQlzql5fBFbuehcCreKTucH22MNqppMfisM/Ffl2HvPdcJyIDu6aRWwuNGWA
i545rNxnBa6M2Iqu6Li8jyqPTY9ZBFFMiQZ/tYoR3GX6+es2d8jJZOQ697papNS2h+rbqMjAVlqJ
Rpt0HxxkJr55PoEGjklBuD++ucbKfmZnm7kiMMDQ8UdRMYj3GJAH+3XGrW2ZiaM5tlcc0sNRzsHK
vTH0ordQN1fIydQXnjhGARRiB4y/dXa2ZPPpUC8KsH2Uzs7i90MbxbxLHxhOcoD7BANv0qufrVWR
sGrV1DlYs9uCXL0bl5qGeqeQdNQCetqy5zzpDDG5FRUDcx6/DyIjqtNEYSpXVEDgkkDMKRTXVehh
xfdPfv4Fr0Jx3u+O7/U8aV8DXU9vNkJ9COu51N1xd9/jrdHHEa4QuzjL+1wxJ1TTqwty8NM97GKJ
Lr+4GcutpvR4utnV0GwQ8SxPvzHE5PL1A/iVS3wWRXQ1zCRYRFv+gwocVCeiT7Um7+YDRi2Dw7DM
EV9Lp0TF1/V0PjkfhUMcamX81d5iWUwINZqadXamkQQrKbysPTrIp4CIIXRpKHoRYDf90l7zZxTO
Qtmm4p06b/QABousKc+BsZJTF39Jqaaq/7Pz9Y47nZ01oFyTJYk6J4d7Lf3PV5NAcg6Ms3JyqSWn
MmZC1uliTzSzoO1mMzPKVrqwVHahFetQGoiJCL6mlOh2JaZ0FrH61F45JeZWCu9NdSPHj9jsaw5C
8Ma5swNeCTSPi3cgerPI/MccSabrrGJJ+UGGAEpsIntBSXVaLYERNWXZBeR/gywYJII1B3jkRrL4
14CbdkfJ9q4wqrQqctt8Q+SGyQ68nWsbvbMWuMa71zZIL4zFmB6nv4P0OiCncyypnqrojYcR+nzX
P8IzZpcbMZBg/eMYQxRRYvH3ijobT8wT4FTuWXuRX1E/xbtUAw4p3exu2feHw8k/m2xL/fTta+J7
G+weaLZFb8K0bkAy/MxxOGdqJfPafYLxcMbLJRf0vB2QAm9lFdLtFzSUlecKQzOjKhgl78RiVcbc
pmr0aiws0TP0hF4ogr5QViLyzgLm7dtyhBhmULJHl6lXQNg7rXQP6BwG0ES4sVXR5BJbn/RN4ciQ
4BMfPMVTymDF0ZlZmmiQ/cfqXw9LJ/7f7tqyST43oUYZE4YulJj/jhelgnu5c9jXGUuiVG1u/z0m
Mx+MLR2fRiWZkqsV+l3CLtKYJr3fQLwjFj847eu6B9ysFhE3pmmhJdO8N0ZM5pAE2DVpjGEr1yLH
6OG9WZQyAarrWuEMYSRO9+eXnXudUG8FxXo/c4a6Jro76i1MKxwyiY7hN+s1KekBQ2dKx6fzGOt+
Uy0xcgjFVgyTtoF/8rBtvcWX+6MBJYq1/n6zMhRVc5ckKnFLkfxpPQHUhdpQu7GkQo0swp2Hpug1
Jke31bzldkhvDaj/KdNWJOUwJsT6Ey9R6d9SLurY0WeN87jc7SH1ceBcmI0e/aqqD7IS8cD6+lkA
Il5kSiUKvbtXa29qBXNOwUtt8RbLiI1n1ri23SFgOpVlDN1dxpiuAtdRWZkGBmfykZ6nZFiVANu5
PkSXx1w1lQ2C+mQFAK2PPxq5JJUBV39a+5lNib39xCoadylwbWR/K9tEvCXgMeAHEtqQblVCciiB
3tDZnrJYV0EoS/etxeF149UqAVME5RnoJTqq2AFQIi12HcJGHbVXjNSDT26P8BCbfGGzSUWkRG43
PVn4Z6JabwvgVz0mrWAtOHqMIVe6A5STAoJwVHcFU+zG9UElzvwVYqUYYsF516cPZJh7mAmhtGoV
1Z5PAqlCRZhTceNXAxWmCuINMLpjLSUNR+l3np0mEDygc2VL6EijhsN+cbaqTopF9+eFPdWIAbYQ
gjsm8fwGU9gTfXa1h39a5mL46hrfPtnNHcLpk7QAZnn+2YjXURpsTpwn0LayR1/h/yA9ZGC5uALT
YsQcrgHE+3CjgLktsKlXrxaoc66SDoDRpzKwvLnSlcIOdXY8ojhuBYy9SWX8y5AOUCufVT6t13Mu
W1Pd6WyrIJWTASgEkhNvtCkDwE97QzjctYtebJZz7xQSjBdJJuVE/dfrTmdpG6Z6UmaGgR8x/Ig7
HVOR14bUGLVOyI+fzQTNQy0QEJM6Advm8wDYccEyTWS1ONXSYpLXlC4k46vS9zOLFWrO2PKq49FS
PLFNAtL8fdHIhqRqmMMuKhFbxoA8SFsJ58hh0RbK0KbopoQMZKQDksEkVXhG1AsltLzXcW1KQOz3
qeTh1/OrKk3hBhSgZ/Njp4RZjIamAxnD27rW892DIWXXK5uSYtjMR8kdK4Qgx2nPrf88dwI4ouGF
qIRyVor3qMjmfWmIINtOGmvzsOXDy9OpdgFJLn8sL7b0vuMJChUqtsw34mfUlupMdab4jdM7OFB2
FA0w329ffnlBGnZxtN3c4/k4NUthly7uFZupY6sd1NPBlgRlbbW81H8e5cr271GtPRo8BFGoTC48
1ovo5E2OIpLnkGHvqYjQFlPazGL/U8YoHG8XZr9tBvAOhIFKdcDr7CTKSG6/b8Nxjb+7QY5JxYPo
SXWY3afyu6vbevIucKdhYihcjIVcs5/F6Uak2uMHfWsuMmDN0AzJrWG3OvUGXjiBnhB2GkDYfCAt
aKf0+PPttK+Uwc41h7H+zZjtyNl0sIpc2m+cjmP48s1kHY15HVdeky0FQcV71dUTXy2LgXT11Bt6
FQOIX4EA+UKV9wkpmZqIR9DGq1QDkRX50jv2S10V+Y6jQ1H5GOPCMzNwB79hFkJA8LbiCFwAbgNg
VZvE9AA7mNuCP6rf8Eey8A/JtpVEdskcshpYhdiocAd0NjgYDN9KQeoj0VkH2BOY4rGKdNO8P1An
AHXdpzv8Py3HFn4WMkHGXNZ+gRihQWX8Vfrr/aaaCTUMWsIwyIhUPe2BgfRmbCtecAtbBa0rcr8f
k1W+cgQFFwmTCTqsYElKrAx05nZwLLN7AnZ9xsNefHJ7b8V03DFKuEzEHh8QMDA/0F4aE3XkDRvP
88kRpL8NLpkUuDAouBr8yYGn/8Yyezmu66iZt31hAeFXmV2ciRcwXlknUITYYX9VB9G5BJM78oJA
J+44RWkjYUQEHXBUu50lXYNKGKh7WFtLWp+4oeVo20IOtjZGdv1wlMRQxq5EL8xZL/7pU+qwogAs
yXAfL9794g3oudY6uhZHXODnDS6vLpW2tEeHSR+m58/us1sYP4x5oDP5FroE//PNWADfNoHy9cOD
jnggzRB8gs/Ln+fV4Ype5Kmg518pydzGQ6hmCF+jy8dx+jt5YtIBvigOPYkd1grB/PRjlb878eOg
6YMhGK0hnlCGs+QBdQjXehM0vLHSbo9tCkMxL7ork7liuliTUV74IUoXmF2Syzh+JcqXJaXd0GwJ
MUY1yfv2vTMhprguK+qkVNV5VZIZWpxNTJH4PTcmWBKjnSGlHeB1Z/3oWRQ1Wj3bNZH4jrPOkRbO
PsbzuUwbXO6qmKSmL54zc7G78Y1zmBjdBLspQsmwZIZ3RSnf6mEgE+yKq0Gf+dP7Knvni1/4H9IT
sjjFQy5rO4VatiNYwvJafhgVxhtR0vt5VI9EENDi1L7YVRMUrUb1uoq/eW/bjq4oePv0lZd7DpJe
YiBF9/Ftsile7BdRMuiM1VAQi8GyCovwL2ACqQbj51EYg0LD/49epeHXsHsl84AccRvi5T+zRV3V
GIUEvWG8pxJXeRWbPs+BjZDijZhw8KPIc2JvPq3auJYPuCFJGbVK2VHOK4Pm4gq8RLE5pbvRo2iT
HSc9VpRH+bRQhifGtjMWBPWLigjEhflsgzfF8R3ZNwcHI6him5HbMOttX92zqJlOTYMMwSjyTnhV
wnW9PsIONy2grnL0ZW256g1YMzwuMK9rUifdQ32FY4osYrZ2uQfYdEukTzGluo0VxJw4KXKCbQXl
aoB8gB89V94Ev+ycrWaGzU7/Kh/rxnn3BjO1cnVFfl6ovJiW81sDBevJbGx0iPO3P4U3wfli5uk0
jTObhpkCPpfcZyuGRTINhVX2JnRKtdNLeU/kYWrlspIwybUT76q2GFgCGqa9uPhRQ8RMl0HNvjQH
a/fIorqMs8/Egz3LXVq1DxZrN7KLdjCEWTo9D7e14yEdSBwWrK+LOPgFqCiORgB3Ex9MbaPFHywI
uEYPJQas8U3of2v0bipBNG/gD3ZJrFMP/tSOuBiMhogzlETIb/3b8gFY6US3vxoaJpbilsUNcypo
zhfP3ylV43WYiwW/U/raicIl/35zBbj9JIYgryvIcV3ZITFF2K4dUQIl7yJ7UxpflaXQjvWfeNWg
momkxIe9zD/WvbCU2mqT+EWqfXFF/J4dkLRTOYX0sX6fSC9L6oAY/Newzib1MeEcHg8bLuflL5/t
hobnLzSjEOl1RTCs27pmRYtql7nYGu824daXlVh9ISng7HEos3nXFSQGJIkgs8LsB3LO+RN52Ica
njZD5kUY4Oy7p4mwgqASyIdNaeyFS/lO7I1RiuQdif7TqE08r11yxyj0GDVPCfKNLi+3w4ZHen4K
TolO8TY+1bT28XEZn8mtlv8gTHO//dYlDZ43+6EtT0MoiKgAFHZenNAYsqXIWw0yLl+TnpAztcbz
dJQUlfpjd9QPaKfnqDb0XdaFdXoiGf0rKUYQJfSrpBJPn93PvRaYTQFF/kzq+MLw64LRiNYgW/JE
zMl2lUlQUx+2gYR1l9N3sC/sy4eC/1DqfKndrmpKaeN2lOfUBv2K5mWVAx/y5Zre16zT6U2vSW01
7K3pYfB86ugVRSRH3yBObvS+KfUoyn6n3dJPHKl5KpqtCZYMseMrNNOdHHAn8TM2/zVjWuIzD1PM
Voz6tyIXMsu2hvdSdTWhRXG40pxmlHdIOqM9DYgvJ4y430B0yBi+srsg3LMB68xNIxlgGgxDPFr1
Q6YvbShKZO64mtosfRJbLtJE2st22OXVKEI02s/qMWu6Q1OEziI2+GHuLzTQ7sQ4MLDrovvvBDPv
/XV8+xAD4M2iwum2ItKwaQdnYlUjaGj7wQRD34GdOYkOOqI3WeAk/xSY2daFTl9X26c9rJAWYlwm
rW5mCx0iFVW1kIw0CekbLd+HTg7OCVspzfp/0Hkdzbf0Vl9WFYe4M5S9lSKRYTy+xdIU+jRqMZXp
geZLOfTeOInGy5V17PRnMgcrVA1e/sAghrOjPR4sRVNbDsRcHU+cpqiruhdb+n5h52YtweHV7RkB
H3KcsQp8NV1meYHcf8nfjoo16efzvgI8idZ5kDbrgvkHt0zU7oHuc3EdxHJYUfumPJVYgbjIl7cH
BDu35MNGprNkvuuEjdyVJhhC7kSm6ogOOCVLbLvmXuyNl0MfN6KmhOjfpQAKuo31+mIJlOra1ZkP
PBQ+Qi7H6UK/jXsrQcQbyrzySBDNu363+UQmDo7rxBdicELEZK+xlrl8iozP30277lWiKp8ovKtq
IS0y4DyElpU9SLUQXIWq7kLfam3UPolHTHh7KL6hlmwTkmYLvOdLqZKEfx43F1mPlv+kn0mR3zjp
cHd9JxM9d3XAzqcdxQLy9WD/XpX/7I9bZXKw1Z0dSALW0ubyUsK5V4VOlY2Fes7KWIU9qXl//b6F
9CkLEUVsGGajxFO/8AJ03V0CutO9bTdYURceWBZnumxc8BbgB8PZfX9Ox1vwjB+LOlceyUBhsjce
8WpOURNnsRG3tKQ6K36869gr+Dw70Bny26Oew8CIjAvLnyOw1y5f3HorOb5zcVpWUd8lTgGRnh1e
qR3W3Tm0BGbNKElD2IHeB49v4eBRtgFXZIrSl4PoT0BR7J9KUahx5JX+7mLCw/U+esxPVPCbkXvb
Q/xKE8kOZ8Vxqv4XNSqGEu/qG/NU8iduKZq6ggCPkAkLqXyl5TngSJhS+ISsvut0uylayyTOWE+U
3F/i2xOI/6I+yxh9akuxVVw+YYcW3FnwW74L1lkHqSFMYOu7hK4TPtZkZNDxVPznYcUU/1z/DCCm
p6umfBTFDfCGzBzDHFxpAYzdvMhDaQxZBHGW+sRvM8xyS8JivSdEhX/12/Wvu7vDVS8h62iG0y7F
GTeje4bX9vbyDvHDE26Fu50IrcSJXIU5oTNBl6TRS80307CypzvF8ZxlBIA2UjDXTM5h/ZIOcYBP
Hd0jfZVpELdWRMkV07y61VFG+KKlGPiN9T/5hoZhSg4hT9B+FCs0SlkxhYZxF5fRfPp0F2wqYLs5
GtLabZ8fylh1KP3pNDS4D/kJYatV4lAi8A3aD9kr2jLfSYu9bjGSRnb3AptGL6/SX0K+4zZOQgeK
8fZ3+KxLV/QW5OfBKVIoDqqAd1ymBTvxadN28HEq0xp1cacTHC0QjHgbDQUPhG+lONU/na//NNYi
4jhIj8k0p4hYdb4voEFMBD52nbgEj15CHLMANJdttlUeByI5C4m9SrAAubVj7y+v00kc5tekFROp
OsToWBtEiYRYJCZ2+7k/x7hqrUEqdHLlxBhJzreXXg9522xMtVHbAdSuHiHGGVo4eb/JXSiooOkD
woRc+/RHOSXsn3o5uZaLDEjZLx83W7BUrGjTT1u+qL2Yq5DsT+WtAy+XNX6V13+5jDCXslSE7anM
tD2cOvynpJ7kflqBF7dxBUc3UNqiZj1zJn2av9AWf+lTzjW6CSG5DZiuK3vnAGFTvOIlBqb9/Jx7
rCeFrm1hEEeV1aFVAnUyyYTaU9rwluhsAyUaLnpFH9AGVnosLvpa9G4sC7qQyqAE6fvSaow5oqF0
sQ9G/ecp5iSepPeDrUzOhwJPTPFQAPVDL/P6bRKFKoN38nn0i4hM7HudYNIjz/SUvbjzB/KVRl2b
23/hr6BE4tUmEV2BcuZi1NzJBiPH/6qUeJLtVVBOICg0AMfZ1LX26FoAdkrv6F7F5bkdUOYZCIGd
mRMOAFFbUFnZhWU83GbUOuGXkii5iw0Dol25CWW981aJpIpasnthS1MCPA6mka+w0SCVV4AJpm2w
2jobSIpzJQ9fMKiFEmfu1dWkwp9BXfC0TdsRDViMp9Lp2flLTSENG5OdWr/OPrqofTLdO3vksEAe
jnu0gAzmTUFml9nCicEXvukJGUSjQhrj+SsBrotzMU/ARKX6+bySHMX5pARmjNjXBg471ffPl2n9
d3gl3h1xmz6tezvV4JJpe2/mrroa4YWcucIS65m0q6FK47eYHNtGb3BmULwQJCaYJoGjRIw+1qHB
QazY8y/sh2oQM+jZ7xyadbZyhkRN3lkqe0FXC1Bcl/eE3b+YvSns+CbalbvAnKml+ETajxrdUNpJ
RMpWb9H+4dhRNstHvT/nlxIgfMWGkzX5V4IU5Upg8Fs75yKf9oX2WmJOMJtboyfdGW+/D5DHoBUq
RnXrc/dIaHtcTF0uPiw0BMPqSM9IzgSgcpLCexcIPtWVaGvjUzchs9td1aYxKsvYDJqnuEt1vo+y
C/D1HTOQtj0W0HoYgjoVuZKTyc6L2/0oCBqYC/s9ezb+kng4zxTflQkD70WL77fQtGAWOEhQ7qCU
rIRn4BbtU+5VgbDlfziaGfgZ+Q1jgZuCM/i9RDE6mYDF9RxRdeIeIvW8riER37Pu5c1b17HmPGWp
rD2KXFx3A77TwFk36gXIBFZ3FiqnF/9Mfp5jflTWwCHeObE7m2X85uamloPpgnIlMNhcHfW27k9y
7me9sYDJ1J2VRCtDUmchZr4rdf+ek8tq7xX0+JkT90p1PIXBkYA6SayqEyNFzqh6r46dHOtyRCQ5
xWBfZDLRHcweQtp4k2Qnx93vqi/Z2Jzll43LVHuureDnbZkJCSiIyUcjyz6BuOGNUP3RH3Jnbu57
yTx3ydiDKIxUEjscD+6b9pGdpYKwlOIaPIKtqAvHMUW2DfvMoNwLtW0oUioQyLJZHUzWUHOhj8PU
GHl3iv1GYbsRFfEwiLeiIsLDgEBMOVtpi8ckh+gCZNAArJARu7CxgBBk6kICPuo+EKo3RYsnYMgJ
j2XjO8rc8oahBgIaXh6eHGkajajEFqaBPgTpL4Bc6sGOhiDwGVb+SUIz2P6mFJ3eQfS0uCmjG+w0
Fir6VczA6b7k5v3hhpIAnOfyOSJ607z2N7WAVIdiSDi7WvVg30+Edulauf8Aio6pvOSxJHkkvJfo
9X/wJEbBQ0sHh3nR1+cYDsThAXmgJgEDdhiHMFiWome0jwl//DFijHiuphTntg3QMP/F8qhR1Q+g
sjO+zQr0rFTFZVmIW/d06DFgtNxNWkO8TlimAURmDjsA1O1rMK4iuntqOPQYToT7izdsgQ+Ltj2o
2+Qkw/Nygscg5bgXMerBG3OBUBSjXQAZXu8euGEkVIziJog8MwOsf4M3S3mltF0/wdS+SMIZGxz9
7BAlItWUvjfemtm4k6Ce18FeAt4TADDYrF/cvm20CU9OrkYozFs3pkYoIrKovg6FkouNIHqaMa9b
+ue1JfN/1tmdwnSuVCb9yGkEz0thCvMDsl480MIAXyLe/IIAvvprgmMIf+mpeagAv5d5rgrw6l9+
Mj6LNDK06VyCUQH+eSpak+uwiqdG453+pI+r8tw1Ux4BnnBPPLQZNWGv4/iwZYPcP4lsUzr+a99G
VaSFyB99Tu/vTpYrWkQcbQ4t2vLuJGrmodwP2GRoQb6gU2q4iO50edMnznVQ7BhfQZ6DVUQ+9Tol
v+SHtI1Sw7irwb7hkLfqaSdW515R8TlwiQ6eSsqEXeeYIavPfeJkRNE5uNLYXJcENGFf6fRPjr5h
T7WtG490Y4bOU0bVIr8xUD5LKv1RloPkoo0qoKWPAwKP9glpPylEHkZYcTpBD5U56j86CVPqTT9V
quEmHVpe3Bkv/brVmKPWXTZFeae5d8ijLADbS8dVeR1URtyKHFVP6u2ReB9qJJr+qR+57jRJsFtW
Q13hc7f+ynltXhSsgIsLIFhR1lc1Nxq3pEy8q8aDsrgrFEbqq8LF1QHPnUdNnFBPH6pQOB+CNcHr
fOhRxvjKmtCP532HnYnfujW8G00KvB0XQfDa6OgpDi3iNPRC0mFErX55vuvTAv3DPrtXqhlzvfUv
dGSWZ2AJY1n78VXyfazHrM0M9TQfiOaKJkle7XIPn4lXLQ/t5wCLLX0ByCpGXWzV4U+QqFhzxR4L
PXTH/Z9ohQ8i2EFHafWZwkM2tFdEhpzYCf2MmW3k3h8wF7VE4mnbvo8Bp0DQwLRdMnr4/a7wOIhY
kfwYRfBCiUbVs8OYosCylyXecL2dztohmaBVl1Oy4ojYqQbP1qfL7ljHfbHYdp2dYP3waSc20ZLx
b0rYUtIhXgcHnt6qcrYTcaFK5HrP6SGxVNlBY142CWpKV8kvYs8oKXV8/5wb/J4qq/8JrTSai+ca
tTa8HWROZNgpVflTmxTs/RkGELhys2plv/I/s0SxytG9SL7ywMPUFMboZmO0e7vSrqamLsZL1P8h
kV/ArnVxdTWDukVMoPMT76xWr3YNLjrxYhRmsoqDVGZMdfowT5v8UQKV67mcoZIB7YjF1K4J7sDZ
+1fsGn8DpS6H2oAGnqYVX59vRL1aCR5oKD/MQk4/NKuU1fbr5IqwbpiCmFcqNEc3cq6kFx9QRIY8
0wiaFQpwuBhRxZ8+hoAhbLXP2ti9fWeq+Fz5DnESSuhtyOGhzC4vVEf6ccg/oe+BIIoejpP8khBC
QG1RcnA3kGEXhvmAXQtIdcIFdY1vR0PKMO3++96zckFDBWjQUcnwjSFm1g2fSg1/DRBJ0vNTf0yc
8Md9xgG8BjKpCr3G2lFjuYZIqUxohzkzECYtbHFpQUZF/tcokvo7ScqEWvvYDOwyq7Tbv6y3pWtp
9Kz3rLnXmrgsKOXGYnCj79ZDTzMxJU3PCSqF8ZmBYjNIlT60f/fh/UdlLGRmsgi+Ox3DRvA4kP8s
etWMXG/03v66HAakUt2auUmNu3M6g8pc+J0vHabrtiSLURUQ1Hk+cgiKnHddlrbTrUK0XDfgDbAu
+q92ItKBFf3EEcGXqtunUvhdLMSH1O1I09zojZIoihRUa5mDS7PRGQr6NeCr6rTefQQR4dk8fiA1
BOY36QZYtTJ2olKT20sLS3VsQQq4xjFpbyc8YyNJWpfx3Qei/WEX7K6Hole4kLIT1/sYXUuVS7/B
dCZytVmRUzXUem9VnMnXa91b+iDuiztBAXy84ThwI5+DRifmpO6xyhmZmn55uynIG5gUy4nTNKvz
SMBPP8oHltRCZowrFFvCQh6fL4NmNFHEEbN6rlO0vRiO3Op7eyCwh2s8VnRLigwTTUUR4YHxYKNf
WY3LFTL7hc8cXCTd9548TVDy3/3/aTwHHMjRZNOzPzg7Y/qUPHxaU8cfd3T/ttzLLBXLRiJtqeMM
NGYUu/qW+jshZJaSvUXAHs4S+aI0K+KIvVuHVBhX6LNFuiCqWsFCsMeuPMsMqe5BFu7u0utKL8k/
Lq5G9IIwlfmLuPDGd6lJToeS0cUYvd2QccqWXLAtxjs5uhOmOzst5Qroir2YbTj7EeVhXg3eovNc
6OGJcOgiuEavFsUVnmzq3tH+QFEqzBNfoi+cNatP9J4nVkeFsNVgIVkb8ll9QU1PTXYLVQinPz7S
C1U7dKD75OD8UNjccj9tmdo/I6tAD2k7IBXnGmYvhVFGWDPh77ecyvNT0CVOuzbW5bIjazeaItu1
MYt8tPub15c5E273zj83vkuFitvPYAt5ngBH/SZkT2lSWA2nXMtW1c67BCbe4VYLk1Xwc/8I3GiY
DwGBJvGEIdK9fwR4jgoO/IorqU6m8qnZ0VoVekkzvwYj2U6KJrCHbgxn82Ww/NCVahXNOIl7Y9zL
zOn7DfyknwEzpECXU6HY/witYJmuudAz+O+qseHI6N+SBiCAShLncb/9iyE/vLSi7oblQgL0w3T/
SVAnV4pK7BI9BaGiBChdLldaEHWO/6UgTs3DprjeH77PXKy+J0fWnxwLAXSl6MnRDO9aEkju6xA+
QhQ7MTyHEW7MZiso5HyfzPrcqB5cQ+GZn5HpN27p5/uynS/AQm77X0f9DigLdtZNwlAPmVNjbnQu
TpYsFjNcijDcbAv93BV6hQ1J9onMDmPpBfnLEoHAv6kgojfJHfw2xBtWz5nqraiwC1HD1Q0/FgWu
S7yl/9YvbraTyd6DEeJIvUFG3mT7uTKh9RSB59+Qw2E4Eg9yspD5FRGGPmnJcooKlSCfrhQed8HY
1KUIAz1X7iRSjme/bWf21qSZSGV4hHqOj6dQbOM09SvXw1olcAeFb1gets67cU05NDC7HAF7Pvvp
xrqRvnpZAgO+0RnBnQcf1BzZBCAaPsQg+qLaHNwo6LaOIihGh/xnEu5jbNab9GIbzN63aP1qQai6
V63c6JKpfsAuKdZQF9ZkFSf1G6GuNrzUMATEoASaTo8XZCDvsLrgfk+TqqRgnABhOYRd8ksK42/s
pM91eMobXtMAYslJV/5c6Gd23+gre+WuKZ2VXovhMpglqGlpVwwcvxwKilqm0mEn7Kpm5+KbQa/C
bq/BylHEwKaoZ6OTbe2bek2/Drc7DinlBxRYqgswG7OHMGbz0YBOkNMY0LX1cBNR9J0AaOZEp08r
/z3Ggqsm44pNL92UUORcNoFBO43d59Hs28oCRbd6UrFYMvFj3R5a2HYmaRpxrlN5FXEoY8gqk/nN
fY/b+3gZkOxWd6RSi/CvF+xBbUnXj/iL5P8j8ET19MXHBvabQMeFuEZBA9Yi8NLhRNrwrwuJ9ZIY
4GQxKZxYSswrfWO94vWhDobYPn6P7YoovFsxYO/fCR5vnn8PI3OScHzLUcXA58pOib+FtSrKYECN
EmWUQCvjfoLgjkR6VbGVBTBzmgTUI9Qq4hOb9u9CvPAFhFLwtaZIfDtAAJjYYVsbzKxijUbWalSP
xhblWWu1NrqkjPXEw7ndSiyyzz007c7Sm7YzYvJbngg6gV91/U8wY87aXqtEZwCuhSk8x8fTruZL
E0AJPEXUG3k/InljQxYmdaq54X7OmiRE/6qCK6OeUNbw5LnTmGcYuJ+gMBs2zL6/wGDff75ELuVT
eNNiTZqtjP5vVg0IhzaswCrAqW48hkKDfX0ACucogNcV6Zl/FpCU0gDilOnopFHGet1zSVSsLjPs
kOYWSySJWUruj237BkeOcW0DEk3CE/Ix7qiI0ttrqXaTaxYvWm1dcojwwPYOUHxDGq0gbL0VcGNt
kmnkCHbxRNDZYzH26d+aHJJcGmnFaLa+e4+Jcc0gwfygohmPCyVn/sc6S38Z+MBM1OKiHTfJtWEM
RXEV+eErD5ZxZd0BWuQwyOCpd1NEL1znsw+34u0dpaufGql14D0MEzefAbW3ZqugyqAvv+yOIDbJ
GFEo07NoeMEH+tO6hEKgT+tYtNTVr3oFM0D7orWGAspa6r3yb+o9rAPkgrB90pjOyx++ey1Jt4Sq
Rd8QjBWZ6uXIMzsPgo6CwD4PdueAO8GshDEQFyO15FDIBPOmPgAmjBf+JnQkgJKaHxCb1FrZmo4/
pS27URq2skRdCa7Cy8BMRXVIWNRVLJiUzrSCNJv2cbRIPnwIC9jdpPfXowkhscqJvIfayHZ8QmqU
pBYFIP97qNq78HJ3kyhQUDSaQl1EtxWYGSzTzR89XvRlm+SvO4R18gjnPWEF122cDI5TCtN6/O82
6p3MvV1mPDkb+vD4MOrVJv3VSlqEdUZUBc6/MXOmkkUCzSEl6XMnQ99bA8m5F0IQRuwZBCDrbPQA
dH9cjD3gFjCxvhU+EckuQN/sv/Os7Iyge3o6yz8H7Oes64Z4uBwTOvsytfQynmp0TCgAVVCbJc1s
PLiaSQ4QtnjWhcpqjhDL/r+cSSd1V8YQJ45wQMiCxVJSP5kkhxNvy07E7NGIMlt15hPVv+Rtj8xG
RJulxoU7nEw5Mmo79jb/8+jJzdfXrPZErMfL6SuM+4Wy3dKPlHdTt6aAufMehW2kmirtL9CLCt2t
6brK0Jus5WqJJOq6JqbUdRivTSKqJ9BMEYrRvmhVwuBytJHGuIrY41GMFOs3iQEChcWwlCf8Hp5a
TNTwMMqZKWvh3gbK7QW+vmg6hzTXSP3TcM8OhPY0AKXize8PBt3ZfWPtxzkj8qRAnJKR+VHFK0S/
cgLSeaLR4yOs3eakz+7//DTDW+yOXQUcCy0AoDzWKGXpNEHFx3ulHwzXug7PzrjVqD797Vc6wGVX
XuotCJ3QYQG6Zqt28i+tnYbbct/+BhLNe+CxPiUAp88l6HUKgi1473zgBon9HD5R9Z7pdzy8clvl
+earL1d3WzTdnsk7WaF/6jpO9guFPDEcQeKY5DmWbQmdF66fXy9ylDw3G3Cb6vwWj9XtR3wqIrkZ
J5fDPv6ti8dBd44Q4BZpzKcaxaiqD/U4+6dE8QJzgYmGVLbwPtTRe9sYulYs0T9EZfpn+e8zqRlh
WXfHMqY94j8Y8rUjdzLq3a3EaPU3zplocTJGMRc3yLyy7GokXY5EVV0QIJGR6YaU1th4we5b9xRq
gP3mY3QuTnC/fOvSaEW7q7GaviIrPw0WF8v1EFumAZr+GLcZPyLwLF6ZhROHZDl/AutfDeqNdaL9
KEuGxxcRffZ6Wo4lIxXmcx5EmFhU5kU6iMzsMhab4XSt6+i2YrOWsk4KxdClEh9kvdEHUFTVseNZ
SH+RYaVFsB4ptOGyVh1owXYcx3/5ee12cwAy7J2IuzeP8gmxb/Zx2mWE0IoN8SXb0poZsXo5c3J4
U38I2kBzBObP+zrAYWWorZTV5zOYozgzZYf0j9KzTnylQ4Fl7COkrua5RIsBBmBL1l0mCylFzUH4
Rg8XNt72c2XoVbJH7nnMuK7FmvoCv2lx81MZ4PslghLHuiPtGQtCQFkEQ90kpM0DhcvVmhuFAB/q
QkldVJw6gPMuS3oGpn6HXR9zYEPZ2oSBPqaG1auMwIzrncR2DiBtH9uCiY6CdpYk/bT2bVwo0Mqv
bwlaohRUnpMsW0Kou2OCwFicQCcnrZaabQzcVd1CPlFlJrJBdrFPXYL6u8KiAJnZW+Kd9n5LYy99
szRV8m6cb8ecps94C4JdxLCDJf6q+kSxr7Y3zt14UuZA2YdSm4AC4jsna/HgUMXIMFW2/b/YqUqR
lp514HPcU7aZdnCCUpgijvLSClZFrG5ABt+iyu1ybKLnd8aR39oeGGMGy7e+cfMFG1yXMHleYu76
OHnh5Zj0+XXCiiPLzGE6AqSrYrGQlyORRUtsFM9tWvUetBRAU+ruQaY2SP+gxt4tIdmdl+DpUtcI
8rPR/hqMMofpUOSDdMANTXU5l6P3E+2J2LzVILHMXyvEyS69Hjn74ZOhOZNnh90JbOGonk0lQ41E
GXqzuKY+WCLgXkm4TOkfAUA8eVKDHiUpKwm/SrLIbaDrtq86BVnkZuYrgteJ6vg7Bo7h0U/XfDOf
DPLGqx8CkllOybE3s21iVBJr+uzkO36+fePee4LL/5KPQ0KhBVTtAD5VakLCJ2ubapvf+JVmnSed
z1nobEVzsgY6Haqhyzj8HwagRLXZQXD/8ajCQ6YOaxwMzUMN9DqVfOS+MDNNI/kUZ2gDcNlbZEJH
fQFgRMjPe1GcsSGiJ9wPfyZGAL7yeBuD7qKwq0PJ2fQM2s4WnDC2raArnqcTs/8zvNsSBJgMg+il
7s0NOym5ka1Hfs1EzsY7pRQN3mJDL4DuKIG/SrdF3YwVdZcIoGhD42Kxwu/KDbcGjxNS46Ajd7Uv
8p6fNHat2KKP5xXtWb9K02jrbrV4/cUl1GMp9e7TPYHR3ETKjJrElqTpMeZ0M+NvPjPKepEAAHo1
jnZ7IF54p7dZ+LFLTFEyYCiPk1fl9gDV1cZPWOoVr3zBiVx/KpoYNnqDCMktrnrSFxnXlAtZuZJL
usDekHvX0zFydrwEdVh85Jnst+E1WN+VvYJ/eygo0cy8yFTFru04R4peLzOwk2AfGI2lv7gi1WXp
XFJFa7uAkPFfJCDxIH9my1eBQosUHznyjxaSkfABJdhT62SBgyCtyTKDxeElkQgPNw/Aj7Od0QWr
qGwQOa1GEolp9znidI/MRjkGs51HczwrSltEVBmA4bawqPhPv/tS/AfMGUW1LvD1haV8rSmP5aVK
FA7vjVc9b1g33sjRpZYjwMOmbOIqv/n2p/8nvMz2H2AFT9kQRSiPsUosB0zQsXZwBSnLITaIlbX9
1sknjvIVXgBjUkTswqs9ueBN/wknXbt1Q1o1GaHdZi6MnzPo9BX26AbjLepPMHgx0xbfH0puY3fO
VJMnF5U81GuROVBacwbWTTecXRphcBOcqIUDJZUUQfPhS2ahKwp2ZWlzqTUNU18VnGmiV4NwDSOT
XNOLfbOE+mw9ajBP2UT61WZYrt2kGG+/XKfDm4/1KUujDmnnWFdsR5RkIoqtB0ejJXi4Hhc6tRHY
2uNRd3hv1B4G3ANMRbagIxuvlKhjc+YZpipsRQtg0Sjuo1tzJLPEbSZbTsaISEC2NXhBywUsbI2b
zdhzteYO+O8r+tVa8Km/5/qtqSSgkEz+A/W9h/b4eaWOvQKdFQZUTAGvIs540gVwH2O8kkgraMJj
Mek8//mWp36h82B+M0bk/+OEO+G21U8sUrZHyEH4ElukCu5PJ138dOxF5c3g2gfezNz8W8zlXqPD
aGP0HtJxzzNo+4G+zORD2WA3029heGZnWb5MoVvHfMtIB36lYDh4MoHWuvmD9P3B+gdYXplD2dMi
kcfh8MeNWZpcv+sL/og0VuztXQZlhd4BfWTlv/xM6b63+QhgVkSj9zoWg0Cv0nqTdfWmOJaNog09
8hWioPIAptZ3R27+BBWrluvzzcy4duJo+Nc4ClN9s3OQA4GGE3hsgJpBdyzgQwJsuvpQYmmI02f5
ZBFCYWjnyF/Ag6QAbiAInSjVbHyepiv/j3RRmUGdGTcnkmvJMxN9kik+7n+TM1Eh0OiVjIxW5AqH
P3wCbgqXFoJbSTDZrgVIMyXdp9dhszcvIEkzTpBw+TS9mlWSCKmsSjm5O/kpN4FBQrRc22Pvr9eO
fqpFVxaW7PLRDL5RBnFGcd2iFpC4C3DJ4F7IrVmo9Poeh3eaUOQN9boBQmbR462WzpkbbWgI59Nu
51N1Zmq1TQC8r26+OOkz12vLVfZKM6/X5lnJdJWhzH2BDQ1ZD0ZnxuQxDxcbvsLSAEuiXPbD/EE4
11nhQB8CqhXnSjhKLUUdZjsvbGl475VGZc9N6Ynvx4AbuBstfTnKcsS0bWP1MeaUOWvW+rLvI+Z4
Tb7qw5zXd/am7nr6Km39voYeTE8gtH2iVmdOx54Bj1/vE2/+agZLcZBEFsDzerHVPDUoLbof2gRj
C8AmGFRgIAo28e8SBkrQCsDQ6xknZJ8TqDf14arTYYZIl0u2JXzo5ni93adcdbBfLpLFqOSVmTRH
0EE7695c9IRevO6v59CYNUxdmhU0eHrD4Q82xhB7bkddwlVcc5WHi4Cxnhn2NFAg9VekKzvonGdc
slqkOMMe5rfB+HuYvjSSnfGZ0C5K2dMpuzGnrWeagj57fFpeTZmoUpIg/GnzFuhAnesEuAe0/Kvb
SLwIs+LIHqFK6SliV8OVQAhnTXglVX/3dYmo5EaseQLmH/7qAMjsP3lnc3sPxxkoWHjr/bpjYWB8
oEmak/Z/xEEts22iU6UdD8Y4MmW0VThhodLvON+hT3X2aBxQZ6j4qrqOeSfzO98bCefw598LVCp9
1b76dPgyxxJmTgYEZ1PtPwg0h5tlZzZAW+BFdaO4uAGAS3WCeCHZNr3BVU45yjxFItASH5xtmQeN
IROCEo6/GbYukJUPFu4OU936BVEqLvh7QJirwlIcUXI62H4Ps8tRO0gC4NT7IRN70PM4yLj7zcGU
JdlSYRrpKw2hyi2PKHehkzqU/nP+2lFhKL625LRS1LHsVON7v5ata6UKrdnhf1uDFkb1N8QLiBOR
r4SLIFl0ySN0pyOMbV5AjrwxuzmlldORzdalXNH4B/Ai6/dj10V/ukvzStrJfrpiSl6ui1vGErLe
gf13SYiHmbI6ThOdcKTLIyOzMyQ8HM1ZH02yatlkp9wBCLzDp0lviQWKVOf1CdpYzL9iBcOpRrn8
QFybznwVBKIqXS3vYMh9C+r1I7qNrqnp/Q1F7SsZlqYkI9lef4jt6yEH8V+i7GgrlRWxeSL4svW8
msqqlK0/S6V2/xM9WnS8L4T4p3TrjbhQgPma4K0rizGznqNLjO6LmG6fuOJPrzx3Dpc5vbhhaiYa
u+7bGyDCDKYiy1djkY88aT2Fi7KCx1+YmsC8hSImlriJpAG2hFCGvCLr9/QKSoobeTYtmnp7zzo9
hpgZACkwWsmqdvddBn9GqcY3PvbtfrswBwuAt08rXRSTaLUIQ2tBAkpkdzENBe4S0LVVzJUzbmWY
fTOH49JcCs+RYbKJcOQ74/GdXppmZF1AamkafLneWrskgjq5pSAjudglg0wkwkLL1KBC3YOFlBNv
uZcBz3iEhXkD2IR/u6blCXNfH2IWWPMNq9JZ0nYaUa4xj2P1IatJjOOoC8+HKgVLgtEiyB2mNCMh
FqrL/yWJ9OLL6rrF8S7WWL9LrVEES4/GDZJda90LGNsRK6MZB7zSuclJT8MLKpQlWYMXlUK6d41r
Y2+FnoKjwi2oKRDrOMtpOlBy10I2ftqk9hD0jb5ux1TZq+Jrfehb8Cyd3JJI2Swxa0hk9AzR3OGC
ONqMdTaFKzbh8NleIHkTyKEAb38d41rZbOakD6IRwf4S6DpzVmc4hIrLONpI1P5DJFjJDRkwEjl4
vL/Ylz1aMdHBHU3YNXw4wqo0GLpN6NnbvnjRnGVAXhRNGwgowMVUW47ige5DoW9JCyNCfSS5jMac
FNuRk8YF2+F7EMtU84Bqz0EvgXX+uf8vXEr+dZOqCkZ7v3dXgkQLwZMbifmn5jmVfK3Y9wOOEW44
IU4hEeE+AugqkMZoBFoqJg07VyIWWc8w9KQBLCUT90iah2Qkjwyl2OuFTCxn+j05bwv1J3D6fhO8
RUZcti4Y6gqHFNaNXEamd/RgRH0bPxvyV0wuL3MyVzBhSRtriuPYZlEoqpnav9K+YaYFHF1zzWwB
3FOrecvgLmtBazM9yhmPUum4jr22qZWxIETgYJOJu5d4T9U81W1b0U4tlHLdDUr8PgJoSa8hgPaV
SZ+XkcfAAQsM0U55kbPg154xRvrx2pmVYSrMjVWz52+oxFy98XGqKsI/ia9uZbYZMAhLL1iwW8wi
UDrwztyNO1Dxxh98r1KQM7sEQcZuSTczq1uPtZNwSs4d1pjXeWhwYrGB/Sx4N3VLrR6g11N8Jod3
VcSV2/MVsDZihYSB2W5gNFhIaduS50TUc7tUZGVfZBRFFn0oFfgsVAOGxdcSYNr2iA+mpiKHBCIg
JUp8DfHacG8+bWc5D0sq+wlSE/tk7F9bs39yFqtt+se1pnsPTjN+XKCSRc2xIQphJSbOWTzsvSgL
Li9Hi62n60KDJTgZdJWuytoyHI5YN0Zz085QmXktbPJxV1dXvLOBZ+/gke4nPSMrzgGEUlUejCdp
DSxd+I/eIz3WOz3Ccl4tiJT3KHGcmOyH9HgLbr1XBQ9eQo32lD6qYIWweu5kgpwOiw1oHu2lyGgn
e3DV+fv8Gq36LE+xy0Trfd6Y12r21zlS127D+hSXeHpX0kqTP1OLNQFU47rGthJBhCNdBQdWdkcb
jlP9XaB7rpbaqd0ROFtoFkVI0T7ZDPFJh+cCajeqdvzalByjqCO1W2nvtrZUXI2b2/ry4TXrLhHE
HPCX8+1tVg3J+e2LM6BY6SpEbgM9hFDyG1C7QbSCK2dfHJEUksnNxulzaEZL+PWohNW+ZTfzfTEP
OuBwd+G5Eoogo+WjUlx+2vo4sH0kQF/w5TbsOOQGxXMpLxqoMZVKsuSj0ejl2ePRrJ70eXQEt7kZ
3FZORvNEFGxPSpQ48T9UOuElbrVe5ReE/RaKIjyv7mBy1SoFGOnLYoi3OQnpQBKY9hTDwQOG98OE
C7xKWBjvOYM0WQewPDJeWMCY/olqvZv2T9cpjA1kYey/65YcoNMQwFugRt7X03dq5xm8dpwgwSoi
bave+Xz5Dnfxdk9pQjsqb/Wto8f69RYjoXTtOMne4DUHZ+jiVdl0Uf0VaQ/IAqK7u64bhMCE/+F6
JndNDnnASlesrKVJ35lipY6o2IgR+K1yQ2MwSfkMVEpD0JvxYoqOBzBkXcus3WARp/MZ0D6GfNVo
HFwNIHazBcZwem+dwuNUlqq+f8rA46vKkWOKzhNpn+YhW85u96cnOoKNs4hXy39rn7MbtopHEq4y
W0rbtLOdr3jECFWuuMuLVsJ1sfE/yI5dOquoJH99eprOQ2zLA6R8M/MBewbSSO5hBdeGcuXN0BLK
V1ZRvwfmLm9om2xx2CmynNHaQ0ah4O3+OW8enHG0EhSTQhJZczXORgtUOsE5NpNnlYFZ7HwlPUek
JVQWHrZ+cUU13jMm9e5BwjXoSTsXQcRTc2P/0xrfupN/5G9vMToiXr4Nriz26H3V0FmZEPo/pIKY
LS9b38E1xM+VnA6rL+TEPpdYvnXZWPlr5THpxTrahNWyzsVdpGkaslR9jYb/6Oe2pjl44k0GYo6h
7JPDk0P0Myk6wuhWYY+xOr0QO9NjIK6UWym0ZiKVdoIUq/bsl6PHnO8p2TkIPlVlyF3ZvqD+6Xts
mwWKGkH2a/4C+W82PZWGvVjZrRbJj1G9Y2g5292Nq9WYofP4d4pV+NRD32qA1obicH00+8VylRlv
G7Owt2N2No4pfy/kUue/lSzC/NitJdsjDtC9pcEoK94Cpe2zTsxG4CIin5sbTTHXTEcSFs2M6AGO
+8mcpwZXaCh7JtWuho6xRbqBRd0HG+4NnmrYUu0ena86XcpPO6eGHLZUpWEAs/4rI/e8X7cX7JMg
P5ijU9XqKFWroyJUN0Aw+UmFql57P6bzOjGhBqG7wufnyBoRkU41fr6QX22B6ucfknirYl4TLPKn
2ij/2pRGep1pdZOOTvVQEVWSP7GfKJwod7ZU18tSiPmds0F95Bmzr4wWbzIXa+cwUZHy+iN4G1gV
BheZ4eX6nQLGGoVjU+r4/kzHnSN0HbmsqVBL57jQeg1e3H/rpkmUsJLlF7XqJ1b55A+5N6Ay7Qvp
HAIOC7KTkGCcF77WYsMcyJ/zRDIRG8JPRIuCsCSjtbetlTKWthSox93mIlQ4nt85Tob8SkohBF+H
o6rNjLzvEjYx34jTOzsyq9PmKyAMvKoEbVLS4hwmxh4AA84t2zG7QJW7sTeQMZ9FGVAmBltRTGlH
uqPkeJr5DDTWAsFpfAPXM8ShACCsg9EdeilcB95MmJBuEPelUcNI/7KDSwXu28raTzJe4a1hEB4j
uRusz/kiCKMd4elQuHAsuRawFsaFrN6NLjNqskJfrkjxzmncBArMQ3sgDRz9v/cmP1UwyHCUOfI5
+H3Iq1RHGlPdYA5+88ZfmRzjQrSH2Wak7/JbFzhKyriYBrz6eU/HNhvrI3vHc4MoiG4CjbKUf1bJ
ItuWr1FFHFGh/OxFXMKfa3zrqNTKiH0O13rfPCKBS04WXZdOWnA4ypKV/Ujr9xW3UZh7QO3x1W9K
xw9rEj9zrSgzDzD0bi1rtsU8s/gkfetvGTfeK4OiPk83Q2PwLtNvJR3Kezp0Mm3t347vbKYmQlCk
eYvqnYeHNT0yggECJTn58NwAz6ZMTPwhPFHaBdRhzvlZ9dOUbP7+I91MJB32JIU7m0JK5vx8s+W4
O0+qdv8AMRddTV8raORZOEU4DOY3IEqNlwVCNpC7zjnFohTAKW75To8mZapsiRiNoRhT2Duq3thG
pg13RtQ2K3na0xnc9/BzPZBf+NSVm/kLf60e4z9mLcAuWxczBqDwz1UXU6QN5XNeBgdcPg7+NcSE
ILYWd1lgCiM/OaA0nEGb23gNIA6Ltn2uW+3x3xUjHahTDnly+1MTrYmFBlk4tnOL5pQDflmsHGGA
+XwR6WBcmrjXWH0t5+19cFiGMAnqPpgduRGWOzQoFm0knCrFQC0olElkBJAwJOctOBlnetF4uFAb
jRJ+7uwWCSjo6g2kcDuvCmZF4pwdrgAFXhyEWfVYV3SZQfU8LsuvMYbu41U8nttmTCEb9Jr3ZBbV
Ey6kc6c0FZ3mQiz0sOoaBs9T1oBLjFP50o9Qv/sBvwrQZ1mHWEV0fvVFJGIpUERrgISEcKGNJB4g
Ne0FbhJUIKwnW68SaQlf+LVCZBPTeXVtLIOvAv0jWFSfvYg2bQzps0bopOzX6apI4Br61QTiEDI0
UJhv98Dt/SdnVhZVdnkUZjVjsC7rNg9t2c+j1gwRB2gKXeWku08ES1PHLmDFpZnoWYU3FIBMpdj5
5OqZHTZcGtJ06XTQ+JR3wRjTQB+ENhPqNVjBeZxrTOo6BtStU44Mb80XB5PSBR7VNrG+yK8LTvKC
IKIkrWgfVkiqjV/SE5um0VoDCy5p51WLU4ZQOTyonNa3YJNNccELiJ2TgorosQle2zfgndRWW5gd
CM95AWzKF31wBYoK4prS+orvSnDiUdx3Dqznt1ekssG6bO313tjbSTaR99vH5q3SESbDpjQfj9FP
ufkdbN9XS89cd2N6oLu/zhTwKXEpmpIjZT2C3kdGTLfa149D027Q5py/Xdt33jfyxWoA9wuvA7eD
2kX6S5+Y+hD2UCBSU/JOt5qY8AEFd1YqJxL7CQxJ+AFy3Wuj3V0WvGeGGDrUSHzZFFgecWnKQmAP
XrVLIDKfbwRSIdqaL+oIFyY+GMvQpvZxxUVgVCLumcAjWRUnK0KAaQA8ajoJ2+qpUW+Se3N143Jl
rCPPK7g008M25xe55UgjvN6amR6k014AWDJOq2Q3qifQd8LlEGEPJynertaW+8blpisIZPD0UQrk
bljyrNpuFO+DK7pYNHkpBuzl1Zz6WSQC5oIQTkV82vhLQ0f4ivb1pY39q2LzObf3R0aoepHY4bzt
GJJ1JvmF+onPsjnU74V7rEugpnn+pOLaMnZGJ8FUVWu3qMa7/0xpKO+cHC6thruw4aZADaSQbT2e
uUk4kt4yHT/9R4dqxVPo34nnZeEMQkci/VXSypp8zO6sM6NrYA5vhM1thDW0xMCUC15y2LLoRaSD
14jcYBp2nwD/9MrHOQBwAo3dZICPHouNO0irg5qelEbvpKSgiWM14pEaGpT11B23m9yTi/jabPLK
Qa6OZubtyILH+Hm1g69xZZvZjfV8+M3jmJC5QO44Gu2B/X42DH3cSTrG/3ome+tYvv/JU8vkL6Ha
1SO80PBIFy0rBbuCyR7xkUbdU0Eu3EeaJc6y3CH11DjxmkSdwUCjYPeMrbxQCF9f63mEv1xZDFkZ
zVrzWi1otEkcSZVGoYnYQKLO3xpmREQ4b8OKMs5Zt5pvpaivz27jWHVc6ptAySBFjkRHD39JYndb
txKpL8T0ZEj7gOkuj7LuBGagxjS0uCsWVCfHYQwOs4t1pNNDsq2wJ23//Km5oL5V8uuVTPZ0gWed
t0azFZ9Sxf/xPv3FukSiuQN1Cj5x2mFOi0ApAt+FgEoDYPBjcTykEC2yWRHW3qYXAoSkInxnRWUX
tMpFf3Jj8ffDCsKr3ZvwPn+qYJR/L6hjBuHxuoKXPB/L0mZLYKYkt/B3qtUvntQCQTejdM4ScHmr
nIGVzIhENqNYoT80Pj+6FNyKkm6M2HyLmy9hROICsDNZvxOyKZKCrfgH8jblOvX52xGo++nMcrzO
DDUnIeVPIZW1cocTWNIHmD8MxUOIRv3pBvlLYRcGMNJsMIkODiq37I2rTQB2+J3BZUQt5ZD2LLom
7ModP4F/HfhTfclJfcqEqpwsyItUdCeqvHyzYhUdFgxUzeyTY5QSO51q44E9W3PXdSrdlbd57IVA
OEtX9ey7i5OPbqlk40divSZcoA36rPWPcLDoknncLrPr2ZjfC05rkfCDhAkMtkR+y7s7BqyDPluE
vjDn63zGSc9PT2V/Ul5FlZF2KoaDeUgocv8c4Mxj1RYIKv9gz2yYA8/Aeyykh4qlQHJVD6/cMx0j
Mh9pyAzZFmzE19CVDelY0GdL3XPgI1xQrg+GkjATnZnrjm3LdGlIFW1P/AY5AHM9shxf5+WEPreA
4OKXZ5q/SXGyWNDhT2qdK3js7GSvWoCO1K4Fo8v2Mgx0C0EhCnmfbfTY5JdfP0mffPPnThyyIrXh
eAT3tzXkzDaoN8S5aVwYZWf9oRb9uxXI/6T8wiKyUpnypNaVNm5I1MDO8DAK5DaEwhLD5Y2cIuiC
TvxWEYbDUlVxmi3ZMSSkOIanYw1mAtwd+6wdRaluWwDtooNHmq7ez1FnO1X1uzKLBivVpgpy6Xpw
7XFUafpiXnG4Eb+u7xBfy2BOWu+cGHnkZhfHAtKOj4yHoO3X+vWJd5xX1WMCNYiYzhmcrqfzz9Y/
p2gTfcX9r65Twl6eFf7u4bJYHh4/HfTNkVvygK6+hFVl5W+Z6aiNWzpP2FTy9nMOMhCL9ZrHiSdB
ptSyflqrQjMPNyI91HXV6dqvFwz1O/x6yNuCtau3DHgVPCV/FY4I0gssIJYnZjxjJK3UiIn7JejB
YTRP1HJcoQNBCgFYveUU3oTOv6y8OJoQX3DO0iW3BgGL4NBxTpBOOWIdqyf3rI03zpSrwtXl9ztV
ogq9H5Hz6mCHYzb9p435C9wYSy4vYHZBJ7RTcfoUhFzxpVIZjnTT7nCYA8g+ne5jpn8f0icudhar
Un++Rn4smLPf+wGvVONCgpOb634faMecuS6kq+Kxr69iO8o8/NgolM8aTJFw+okxP3/M1ZKGl47n
NAEgOi9xDiR/1WAocpFzfCQsq2sC0ZSItw9EYTSh/L4pt8lZdpbIOMM+pHm2q2YnRhvPwCjleMsa
R7hFJwKN7Kev2VNjbydI60ZtJE6Lxpv0sEcA237cITzYtekxdomoVc2XPGyeAEE6JtHpCMyqcd15
hUliA4uEVEAH0WkW3I/7R9hnDKzyWRRgouYzhd9TLnCRwalMvLsUFv1KZlvy9+PBliel9G6K0yqK
lPhspFPtpwBBvEPj59pGNBrCeVMYPpkf28zWDxCakeOogAvcXmTq0ZaP5Cs9KD3hQa1Wni9xgWsl
r0MMioInwavH3gs6+SLRbMT7snmiM+rQeAPQTZ64OmtlF5l7Cc2cssUB//8QUoOZ+COc8ANETYAn
06q3TZSeqPlzOdHNJA4HnIIWHZkRGFz1JyDrzcI/E/80Tsn5waO1sGG5VrDuhxH+XlOKHz0Sl+x8
bm3Y9TdS3APqM4Zw7mAOxG4ELXeyRXFL9a2/cGAjjPgDa1Ktcegz5EHfRpioEbwQWxWoR2JSAPVa
PbGPZydCB/m9hJ/X3iV5o91F5cQpgTaWhZO3Pfvq0dGAcarDvq9ayFYbDB+jSxjUHj0yYiVPDjtr
uhbqECzZ5x5JVpYZlhJ6pf+NhY0fQptayXkpVnnw4f/iD3TuwEpLUCrHqujgmfiDgLciwihvHUVI
+VzW7ZxZVmTMUbIRGIG0gntGvenNVj+s70uqWdhv5E3D8pSGj9rMYIdhMmCVTQYC387Ii3RELubO
qr8qnV+gCa1TXZiG29TiEaUcKtnTVF0yofdngfQTVblw0nNNMgSfe+osgaSJVfPBvQ3NBMWtsQh8
VvEYLpM8z1zRBWZzkvL1ZKbK/c7uMzng/szsPzBYAwerWzxjnyuSCdxfzuDBQKHtoJiWhRAdYibu
7Ma5wcVgtuBdhDBHUrZdpCqdd/fW5sB8nZSANBUfHx9NEwO5CyY61ZR0GR9SM3yUK743PXZvi4c9
q5WPTX1VrhNDS30zsPOzKqguL6oB+HRZ+lsMno+ICuYru6bOqHMFpfWcc7drcWY51qAIcH9/bXjM
u1JeTL11p+9AA2gpSYRapbdO1jlENYif3k1ihBwYjU+K/r54dKiRT3xHIgl2imacHyQdYVPmotqL
OJbW3ZXzuP64l59+geGnDYWUfAhJks42ADtgbnoHMGocObnNTHjq7eaQnmb8M/HYCbAE9ejlBfc2
WnKaFbrf8jWSiZaO6m/skY4VuGXvr3VESZWKfnFwkPFdwYckfbZmun1s1u+0uDfboRXgv3WRTf6A
aDdDKb06f4ARKmqWo7jF8c4VbnvkUzmvVe8o6aEzFepR999Ll2/8BIESea1JQ3WkMcaMlD84Jlmo
AIyW3NYH+O19F1r+W2OYJU7aC34xbObmjOwF3qWdw+PwFtj1I5ohpXmTrEVzVXqkUWwAyYpkiMHI
ugd+mc2zlBYtHzmtncekpB1lmN9Smm1d1NT2sb9spaA8KX0EA37K81/sJN4c3t+5D4qfX82xDkoB
AY3x4+RP9SKP6HmVACoCNCesTiOGCjWmb5X0JhsWGRUT9Vwnkaz7gSSX5KPKmdevZngmYkWq6GGn
X/4YSJxmhpLccB8A/Yr+CwRHl7O2kML8e6kexdzL0uWSAX38CvzkmbK4zXP6YmkhhI1Z/dDkJHiW
QqlSDOeARXz+Zag62x2VRrIRJWETPONF2l8pHhLHVr3vmeHa9dHG7GdbpoDrgXf9kr2CXBkOZuCD
O7N8eL05kpoqcDVoQn6U3fgDgqkyQ2tvQUg4AybtlfAZgLWGx5I/2LI4X9dbdEidBRLzdgniwmvA
M2fNMmti8PklIL63Q1qT1lnEDeNRxKXiXfAcakpObwX9RCtlw+C2retTo1J5e65ENyIfBz6Qy3JJ
/MWD8t3Iv9kcRiiSOBgGAoXNYNbEZ5Cvn6EfYICPyhoQoLKVnFvsniUHyGsPbZTE8WvGs5f+qDjL
r/ZiR2xrOvQ632Q1UJXKItMlfgv7NkzrMogi3GEDNPmjVEZdsz7/y7cMz/dgFYcFmLAFwy3GPfdH
IPtg0DAY6CKMXR4kKDaspo5CZx9+QRxftV9GbPjE2G/2eblvahMAHYzi7YRH6+dlivQeWW+uknwR
u3sggTynqrE9cqjvVwmnz6xYnDuR9tFLXoIJvouPQDYMFbO3H/sWmVBL12e3u82A2uz9/8Sqfxxu
LtvxzK9N0yQoWkIFusqNIu1IU48mjCATBokIvgLZlBuV1wjfJ2PYBeoWvS49u7MdSCnkgoKkGW3m
8uRjSoec7rbE2s7fO2HYVdrgGhclZrpVUIDrOdF0hw2NPssf8JUJHXShu8kCJbuJvLzyS83+uBKJ
DliivHBMtLq6y6uyR1e8RrUm9EtKkUztyS5bn8LlZFDori8hHX/1mDeoLFkN8JVqQo50Y/2EHdCp
LvKA0IlgEUz1qkX+9N/vg1bOlwhfpwGYLlamJB8vEPMmsKDaqK4D75iybPKjapwauvamnM29f5g/
01wj4SwsV2vHHl900R+lRildI38WcnKJ/m06JIIBg47Q7sic341UQMib5cVSjjPasFevck3zZt8C
8FxZTF1gc82kq/uWZa6Xm5TrLeQCAWHZtPSqfv92gI4cIKYvmpUDPN6i+756AUny6h5sSXEfDa/X
ufc9Y2q2q1kpt4SuLuSllifauCb8DLAUYgKMV2hGWWAQ7zOR6mfF/S318orlLydLb2fpzl8zXSmD
L27PPf94XaTR2mmMw28Wf5nO3F820p5YIw5iBOpliZJrj7UDljfBe4/chQrG6u1wFuv8FSywyqPb
XQjYlsfXgghqT0jEOjHZufqc3WAMldmSTwWypxBDWibcZh4w0ycQ3rF0nACvRB2d4z4UIDrJmTc9
LQpp03GTSTpnx9t6SVh+itZ11e9J20cMGXRa7ebc9rN9N8RlI6ha8hbuAyb5OupD6NgQ863PFWem
/N+hYnizDlnH9UNm8ENDg53DIIYPcoVuREhMRpw9BIk+tzBLc5IT7hM/3fqiv7D+KvdFpqVI3OlM
kkmFXPcw3q+Beoo91gdP8i4VsJ56FZ+ro/LKNWHOBVKtuSkvsrWib/ChEMH92kPlc5uq4C3EeGjE
JGdHlTN2aFf8E8UaRcB17BcJED+iag+QHOOz/sfWMyUP8EmDMq7ujgP7cZNDq/UmEyhe78HJyh57
gPJWA2i7jTNyhY/I4f3EDfb/jaZhHsF/VcpsTsufcqmyt/kqPYcPymSPzqVBiJhioF71THaiOvlh
+AfHeYYzSFgFYFbMGCCJrZl6qC2jSSmkY+BEJaT3ciemYHxVelwLgQCL8wCQ+EYC5Wy6FUoqAc1m
Z1t6VuU7SAgo7Q8obTc9zBcpzo7j2HlprnuXP9GdqTzL8d/jzzPbYaRl8wDnkdS4IoqUacLP3FCI
y5KCBSOzGR+iKUJ8sM9e+5TYAVajWQt3IspeF6t4yCLbed3kpqh/fX7C+KtbWm1WIgyGuHlTgG3Q
DlX7qbvhtpN5fI2MKhZ91cUFpxTe1szDVYo7hbFahlh1ryMDNODTKKWA73jCqroaFP0tmZDUng6c
uusIq6JbtacxhWfFg7FEbzebkVElRkSeGKLzlswYSjmCVzyCtNwjs6ZtkGmnho6PsswB7VgtLFXu
0kjYrhC14HmQFZ1ykewgmhuiExl3uWcBZgQ7t2JnHT+XkOoiDnfNYBhgxvUbYqKxWSwWSKWMauWO
vMxwYCvRuEJSm79tJl896BXWNf05kOsVVROu6189VZTbyRkkPd2mPaqgr3OiVi4sy+h+MM1MFM81
gqGjigeJN7jTQJzzyBSXmfQ9Jck6bzst6s5ji9omoERp1JipqzOKama0xwwLwISpPcTezRxc8d+e
BWZxCIIdjOfJxIDNkONaNuF7qtAcaUrd1oeENY2syUzoTvoxDn+VL2zrKEO+TTCtFAhCZ0fa1ZGJ
Uvm+HRR7HltHftAEdSx4jPPlClsJVxlutTgf2tc+FHwKQaVne6Xx2WlFfQzW6pZPz25MQlr83nhV
JR/uGLvTAxB1/DPvNKE79YAt2n5UnM9v+ollo5iHGC4eKW4YDR5WZKxx59fS2X0dBZzBcePkoSUm
QdgFlbrVn5gmFKpYMwxWBviwQh9B4rMZkg47Tz5HJ3XmAtg1QqtEl4W1gufc98sRN0ci9mXn7lri
5fwrPFuLytEplara8VPR+e8BmmAs0ma4TTtj7eTm3ACyR1jnINKu1H0IyFxAVLemh+ye+x5PLFct
5bkHCZ5mseTwRjS2lFCPDEIXMD3eeEARr6qKGRIWkDE/WaW9v0n2CvE6F8yL9ktUvSimosc0GpmF
pIMfsLPvATpx1gvIxMnEoJ3wARtF1ssV6Gl0Ry5rmvGpXVIggDw6zg3rvQxOS2vWbXxgCnHU3ANK
C8TBpeftAI15WXX4EBL7njoU218i6ZQsQQ9Xds3ek/bVEXPDRdu5qxSQa/s4XRaM8xdC7srvZG77
a+Q1QYxkcou+KCmkZVwx+WYylmzzQTo37I+eDOPp07zkm9QN5Q5OalLlnXbnBzdrfEoY8rV4LHUm
zeVN5engJ4+ZFbN/N7V3mtbggrmRX8LbJB9/h45bPlWWizvdv2lT8qQerFC/Z4EM4yQkCWxJILiq
KobkbpPuAmTmw8n6ISZrK/xlIPXv/PzT0Wv1HBGn+0oKJKc8oA/TD3UKg6ZOjSNaveiXPhIjZaKJ
WAsNUocwB92vVfepqURviHcHXo8mA1B+SyvAD5xCRBiSQ7swrXPB9NathTmM/IY9EJlIitaXyZWx
nvZr3Nwn2Wn5OIjFvv0rn+xR6urCuW7UxesKgIRdWSuscAycCUWciwqLNdp/LDStKau8kPNOksTs
xQ3sfy5jxeBPeltxVQ38kBmM/pV884cmolG6NBxeO+iKmTzFFhOWQs+OdAt9prvWOycos5Bw1rXf
Wa560OZ/n5uzIK9LoD1w/g5CV7ue/nuwyzBptZUF7OtM5vj2alDEvnsw0ZKjK6StuXsfAs5EOoaF
ioO/E+iv/N0a2r56scNSIFc4jgLc1sBHs6L7JC0n3eK4vhdrA31KaX1L2gTGA/Vn6/GEqDJhlrq+
Vos28K8tmwD/pNPoeIBrHKramWk6HEdCIK5WIot91B5qNqhhHib3KdWvJ7m2BPQltdOz5IG9SBgt
eDNdRjinMhwE4MwBRwgh/wiGwmG+q2cYHuHz8CauoVmjynlnjVJ9WUjZQfCbPlOsyfgzJyuEmAMi
6B2/Y/RXBYetvPZOHDIEoUSurXxJVx32FKKuYYJmaEpukPXNwNQ/02ZfNx8dsy+0Q79QitupanI3
UqEl/Px1oTpaF2x13AGdMyXjE+zVyWA3fDwqOJgrI3pfnrZmvAZ8dtj/SXbBYnZX1Qlnpp+w2uV0
uDLteNLsvCZ3ZzzThcO7Ybz3krKAcgKOTvV+U3w0FHBG6Vn+SE93pWU8v1wgqH9P/gSC1A2LXNK6
aM28BBfUea+idM/dj6RZt3mOeY2Dl9s7nFXt5+5CkqMAQeuAZdNFtDa3nFaEjCrjZ1/Jkj+9Q5Xj
oOLrWJW6d3tudWhKBdF1SFVeMmBrkf2gt/FKwwKSjNgGAjaADVvfM48s5QwuLix1CCjrquiDe15k
ijBEiLmwl+CQgvdp5kQ7kXvdkQX6oNXtdfxNO59wT6PAcV9hjzCt49wEoeEtqFgrdN/ev56FfDDX
EC33TWDyZ5ntN65TEh00RgQbWtg9ODEcpOq3ASjeKjnOW+bDeIzERHnUdKIMhHOQhbjbTcbWjPS+
kqx6K4ryVrgFqSxzu483zSb8ILCieWgqRfdIlDQqekYvhv0Hq9bccuFxYKhan+6wVepfA4CnyL60
h+O/Hogr/maSfny4Ni7olOnX3flvjLN2o8+i350ygooCVKDCMZXCnxxO7QYuCEKe16+JzfMgp3+0
0ayb5V3jJmcXceQF39Jt/pRhErUhYUtnxUlHjp5DgJAWREJSoIyveCx7lardsIjMSorN8l3VZpM9
Tkgk0ZQmtrHOljTegTM5T5KDE5TD09QtQeNc9NwuYP1Ti/a+wOOpnexsJLq0h/2YzGbooCB61/Xw
Cs296BFls6K3iNxsO2b+aOcscGYI2wknU16eE0yxiI/niKvVyGx1ANA+BH5XwufkykoDcFYJTFt2
2o5XiwXZR2gH6Y2Ui1S95L3Mu4tIUmnojoTj0/pol6jnCDyUdW2GFgPVzlq+nsiBzgSPXT7K2bvN
rsrIBJF7zOsV5BO5aP0BQP60WQQD2ReEGidSTWj7UbmhI7cWEVjFgNCkzx9j/0pt6OKTIc00IP+v
XrK6Ry3qWxUtoOZzQHBbUbU0lKh1+j40SM0vOyZ0jrLxh/7Emfeaoax4KKaNg9ZS3xqE2YTpcE8o
Qg9+czquQylNiBx456MZ0p8AFHSFw+QpnGDA4bMx/9J7xzdHKtjJ3dl/i63sDF7CPKTEMjZOXSpw
EOCYw9FUg5SogW5AMuK1bTWbWyUl0FouYfZcX154ut/WHNxd88VEmAs65zDpqY3Ux5SnO+CqYZBh
lU9KEu/w8RXnCvMHViOIWOtzAjSicNMvxIepKTmBQv1Tw19nT3+wvdorV3uTjLgPIavtQMDfgYE4
86H2MIx0C7LRTrGgeghQXYP4F+TV3fXn42RLt/NU9q2IdGMp89JhMeaK8sJxpmU1KyJZo9PdhCZb
45ENaMlYd8zP5pKiwb/26r5PHEMh2R7sqX/OOuh19ZeFr4W05StuZrYXfwHFg2ZwIkBlQnoDmh4B
6eCYtbgl1Dmq0fIZNDHTJBiVTA8W5Oim2Sz7Zgf3DwGCIeANB1vAad+4DyKSVJVPpnzhf3e/wMsW
KU21+SVxCqS/5zq/mO0TNSB5CUVvnIYAPI6mwkzjB7mPIBxsbP76QMwDXzsCWfTZh9/UsjMbbaqC
BvDMGpu4ED4i2bnhh0rePwXnBPWZFHJQV2yjgSkHHye2DCbjU8OE9Ofwiwv2crN1zEaE4zTkMA6o
n+k/Edd4fiKgItaWos11w1tknZSAY6mIafPdSBE8sCKdlBtfT5u0ZkcdZfBHRoqJ/jEj8hDHlkYY
cThef/+DAkFiHsaW1qQG2X3j0sLCwE/Yhr3D/QXUZsAGlVDcgCfDYYSJ3QHRz4MhqtOE/kGuiVOQ
jljPVRpXzRLl9SN0yTk35GrbN5ToYw5M2xE/qD5YdROOzrfFfGEH77JuL0Lacib0n7gXhrBzE851
awo76bCNSQvKcOaj3sOjAoU2DxeizDI/BqVBBwKkE/bCp3w0baTIw0AUtagCbnDUEp5/DpMAk60Z
sk7Jg7p2ICD1E59tILyfc1HmLhVYSYGiGb201c/EZ9iyuAusESeV1qzgCcgn5AAYdeiU+fpieocH
8xJNkomEWIhY4ogsrqfbus0MdoAG5fxpzLDfLrS3EFdSXuBEKmt7nr9CA7Bit73h6L/CFzrNRmHe
tBhJ71LrCPcCXxzJSZr6JbfxRoohwihjEF9E5Be+vNA785Af3cr8FjfLg2Oq4S73NDjQRZHyPR7R
DE0w8FMMmyqMvuKMiHHHRO2I6o51Enr3aI922ov9kqzcOGGHCJPBGsnjrt4FvI0ksuwMYFvZeWOl
hZFpIo1+RgZ5LNImi2ch0ET4fsNr06Wxhc/RitQxNh8F3k5KTBfpVYB0VCE8XvHWdU7JxYXkh0+N
7+mkLZGl3i6PmH298q/zB5y17p06JdmnPqT7ZLNSNuW8T2/AqXb+7e84CK4GRFmDs/xe+38BW9F3
YHD7aonWIgh7G0XBtLUlfjdy+ElTsVv+g1yyZNuALdBrRZ1k8Rzt3YhygsH/z8hb6cok+QUGEYPe
Jc7iOUVszoIWLtjsDNjQAmI9KSlwPe0VYmZFUc6iG8FfeSUR+chR7fW5zAR4hkYBhEcPlET7GfRl
ny1YPzxMhXjebdfK2tzhmpKG0EY97rctrPQx4H3i2nJxLOJlO33ctxKvxSeAvRJJbNwhw/HjwZt5
tBtjTVY3koDOLYqucxKq/USGbahh3IhoY21P/G+BG+VPZz+f4lMqc8gg43t0Qn4642qzbC/ddFYt
gKmypYA/WsOFy8ijApRD+AbBj4pbqSusmgj4/TfiBF2PzqJVVVrn9t2Pxc7lEUEnEuRK2qvOV9YF
gPfVfuAVYcG7LWrkaNO9Evfu/yB5zgWPjLBBkHe/wZji5ECPAtkR/zsZ9RrWjDqcXPn/6GNsWex5
XtVQJ5I/rac/GIL3G4c/Tw13PgZsmeGKGncl4F556c3OWFNUgCnUTPanC5J1NBDjzQxTvcE3y9Yd
7UYZGovvcOC/krV8fZxj/NA99ah7tLbIi/Wi800U6Ao0+A5aW2qycCHTElIAUQnOzmdSc4owZ5v3
1X/kbqGqYsQRUXn0rMox9TlwVutAJ1xQ/3d2LC9EOAfno/yJ1hDbdv/DAP3AbiTto2HtZxejZZ4q
LV9uGS3LlPVrO/N6GwNY5RktD65icEoEBXFih46faYip+Us8hb6FiDmfovXLdDmEBJC6XrerXOT5
2K3xTJwsy5XDAgrJbzi0Wq69E7JgoJFKmDh7OhByKwlFlu80NzX67+XwjuMinHcJbQhQaKOYEhbn
yADYukodOB+1vyChdk3bE4baEkklYTSCpcCajzXRnq9jGGnv0nsh+5Qfl8a4u1MPDV2GepzyMcKa
YN37bgqON5ac56X/hPhHsyMWNID4ATrm0dOi3rE4eZ3hLC15Dt8hE7RM19gwGIRmSkVfiwWRqa3/
zhziT96kjRKBHZXxrCK4pEWlsSsyQ2mIawBP9mTEyCJUWkN/U5UoV5KvPJFJ8ECFzk1iOnFEqA2A
0068WDnaE2tIRY47TxlG9pGzR+LT6mCOxkFc5zi9wo8zWRJb8HxYR9LwgJNZiho7RiSd13ZDO3OC
8t5UxbIsUZZXjulbfoDkiOOmNUSbEZ+OoGSc/pRKxAj8adHXc/g8vg4zl8BNZfRRYEe1/XNHsKYz
rLj5XR/c8gqEvA0BLvmZfSNL+vDw1RBTIg7flRDfqWjRxskS/nFEAfazlkV4PKDjtmzg1u9fODya
cjfEh+gETmpElu6NYHEVB0yhKLnbC2RBk5hbE/HuTBGKPxgUIFcep1uv/Mq2Y9hy7jTJtzrVdtAI
1F398jQysZClqh2W0OgVjb24EGw/OhSXZ0MBuIPPPWdbeTjoi2JziOevjDyX6fud7bUwetKMp1Fk
XyPmJASmM1U0nZTAdFt6PpwQMkChXYyHziJSp3VLj6OSboHdAV3iVVgBXn+6LI3987Uvz6Uuyhlk
73sAWE1iNjoctgIAYBXsOo+bJssEjykftmq+KUi8qYXU8NDp9sE4SwkJIDBkq0bA+2zehtM3ZnV4
mObl5eAHajCTcUJ76g1qDoFAlHNvqjwE1fASFrA5+QetL70NCwr/xG9wL9/tlttxg9Wzje3IY4++
ruPfji6mRDpdxy0LbzFECo2g+dc37Xm6NXjy1CgfeCBWJF4uZ456YzaIY9gF0D7dFfCpSZRJbxua
bJpU7Vf9pDR1gvgZaebqpvd49oEHj73o4XRAlXjzgBz7hG69EK8akefJ3y+GIbHF1eOF+ZPGSYqq
ePiN/8Q1Jh0pdlPhtjZ9biT57v0P/9fBChxDcYKZV9xwbkdammc3ur1eJ2qfexvPp2Ujc6XpO6iF
rNwsARh85Z8jhNohh1V2Es1F+uixDC2lyRzCnAxYhazDryB7aKuTBz10zGHZO6d7ypr75eeJXi3m
kxz3zCLwvLrikvapeIPUh7+bGXDIEKrtrXUDb01BIv+zPDHyziZTPhoaqy/ZR4mEsfh2V7jGu7HS
P5xP6v6U2VCzALHF0vnCyCK2y98fA2d2c5/TsSB9+aX1NnUHF8bpssKTF4Ln4BiOTsah7W/Q86SJ
PgQAJFaXVKF0Wuyk+VtLDI4MXqTNeSKh/uegqK4OVWGJxiBdRKhVI8lPSryAQRa5q9gsQ6pLHCuc
yYS11bt2R1khYXHaFxFtP8CRg5nG2kMK90q2XtEpPTk318i98DMH4EezDlulQ1sQf1cB30REwv1K
7j7eorQps9son95+pE+AxC+fUdcs9byh56LnYNWxaVfkCIHtwt+EDZ0KQ23RU9C9IimaREgk3mDP
KVr42Ovd3ttEFMtco29eu+dKXFgxNhDNB5puRzTO07zlIZIpV0Hu6aGka5YSZcjgHhOPELLSWUp3
cHSAZXofshWSKFBcTzSiGQfjduJuY6kO8n8hfUFPzgGoYL93kEb4iwYUkuyJu0ZY7ZTSTop80Btl
dBp+pybcnCVd39QnyMEolTDc6QrSE74i+NFkbXasDbsH9CjIdjtWdyFcqGg8h/zKfI+SIj0roR5+
uIWLVxuZsHTO7DEKfuA93TVP44WsZoJQdUGGiYaAqPioFUUnc0tRFdtSHVa8rJDLDxw3P8bOJua0
VzZWEXcURinKskG4ArgGQOADPV1eMmJRT9sbedKcq0AUR10dC0cFHidA0L4rzapnLfvF6xQChi/h
4PvVsy8HTYCyWdZ1TGlwSSBL+l11Br+FBbpNFqAteZfuivRz/orKIAl8qudLhU9HQWgNORDarx2a
eshexd/NokzyRwjmHENSAL+t9W1pEMx5bDPGf3CGpE0wHVwf552OjulUJr23HexeSGB+GeOJNNyL
00VrvM7OIvKPyZMqptKTpegJKRtjmBoJ1V0Bq9jyXevuanMeaUQARTlcOapE8NNByaXGLGdJ5URN
DIu85LPRsWmogvq6ZwX/OicMJ1pBfy+8lwMe06yhc/DP5TH+PbWk6a6S5+zwIbwWA1NZL65DDK+A
d1KRtRsGNK2cOywgGuL5CvZyUl8ZbQpt1tMeEZRfyOijUE4K/KHntK2l/rUjH+HJbQXQjhN69TrM
lBtYSg8GyVLcJNPf63s+VHxLJYje9gZAtMIJCpQCihDIKb7cMfTjnuP0MTk0UZeUAKh7VTDO4RCR
vkCTOJlf5/9gXprzGK3aMMMGbeup7QNNE7/KOrfWGvng2R9rIlW1h94/Gw0hMYwB4hFHbsjwhjyf
N1fvTMQ8/ZKyH1UN+CAdqM0wMsEats3tM2C5VsXYpkKJ+UKpg469f8S3b12TzgTIa0NjkqJzEb9d
3BKrblc1YeRwagBgAtQq++O2MExgKqLdKvJvKFo2esSFax28RWxpF/A2o804BosEMCAhc4ZL43DJ
orq8AG6srJvmF94ewi/nKgrm1eMRl3TYsMrk9jjqCpN2AL4hdclPWIxVhnH+MdpeLk4sj+j1t6ON
/58lkh1FHkHRMF7UGe6cusedb8BTIgLFqXikvJgFULTpjJpM3D31o8lWCIap/WZC7+THbPNkg4KJ
Zxt2JllRVkTvF4GumVZXTwXBjVZN0naxDP1ufxjF6PakDkEzpwsdhVyZsV2qUasly7vft1GObVz/
/+bxyuYJTqdy/zQUxfgsjyBqlRK9NTbU+vh9vFOw4dfrzYqIukGmxDWZ0tUplPpzI34vpc/4wTY3
SrVw7xDpkNYiGsYDNPy7wgSJgiSMpiDB499EOCkviylvTzuWhs9djzicfXw5Q3tCb/IpvnPSDuIW
2zA7k9piuwd7uCzA05fJBABk/ftnSUSqiTpJWUzcqtrcgRVLy3od4zP5GD+535H4YooiYV2MRSJR
JON3elerNtc/fElGjAuEQqwnEfayUaBh3Gw2Yvdll7nyPMBz4UsHTPpmBOEMsDdwZ9WEZRSCUpV3
J0Owcz4p2Q1+fcxzgvo/nXSPrsN2jASKk4rzRDudzGhlEaLgjlHxzAfNf+6ZZjt01l45o/8NTMBf
Wwvh24o75mOQiYRI12zuJOtxUdHAfiBqRT2f2jCDxeuC0Id3L+b/HMwEeV0UpHg1XNRk7eFEA7JM
6e8FMp4iQkzdLVpkwzwv123NvRGOHepCpXtU3qcv4DI6Yws41fqBbOl+FDkeG+a0mBdpgjzkGOXx
9+wAaKEB8RPW+ykLxwHHipo6RM8VvLOHHBCrXSVfh6Efi+H7tJldas/LGjuAn0w3nH523cTrEjd6
FHuJxpbywfRn8xg6/NvEdjK7awDQUfNcg/aj2DoyVTALjoWaap5eociKR64/qf7JzAWOFgZYFyH4
mgBes8dfGEL/hZiM7j+ak+E7op5M4cA1D6uOM28IXoK1Uj/XLBb3AqooXyW4r6QWwAdtRJftRpLe
AtB2tgnAv9tz2ZgaAD9YEMzq7RqS/spFWUERlZhsOiMUViSwvECzNGKZB4rALje/Rm2Sdf2mewfU
pxIX8GB16yFW05WrMvBZdIirr5wYCIZRZxD67YYLMANXhHzHkGDA63OiDrivm+NiwEXiM21z2TgB
pGKIrZj2aq91ETk6d4ScvuQH3ApknRm/gvrmJYf7J6ENbinqP3gORoEtk1nEr8i10nUq79fTrtGp
umA5AiZLKenTKDt2WrVWoJKUk4B58AYERmqPuXtaFesEmBi066n+wu05a4S4uCX1YdT51taw1O1+
qV0rWjzz7qKdKnBo5geP6ZnkoR0e/JCSZFrIELqAJQpB0dizjEuExMKyvw/M6nDgcIAcbMY/uUE+
fSYUkgxFdkLl/ocBn80uBTI0M2bfkKpYVWhFXVwL36NjhZu6M+Kre4p8Se9OrprgOIOUr47Ol1Az
TY35VgRbcQpltVfQO2WLO8DN19S+SHHJopkEP4r9k0YUsyOJtFMoajX2O5xDii5bUgM6O6HTDfWY
sedUVb+jW2t/4ubL+rZsDjgv6EHeiUBqX9iVKEUv38CzqNout9oU0/hFJmf/+SPBHV7k+2jkITab
3hNaTgwI4B14/MZpreNg7vLH4xAIdgzt1iKkhNf3SagqOQaqFn8Aggyk7ds2EpSU5sLyvEUaCbzJ
XI7mmhl155u9XGQ79r43iMg5TZ0yWMbVIit9RoHsNok6lvVrGm5+Da+Hwsy8K5uwKc7bPOYUCbBi
1Y0AsJfh/X+/r+gFsxBUBQywfzzbKDEIQoRUfNwhqFZw2NZ76yf/4ymDj5HmiAZnxR5qnww2Vu6t
9Y3hPVlNwZ0qaIs9lDLP/qRD+k03WxdG+4pYy8KrwEtcwIZPunbELbfwjXotosocj7WvZLoPacEV
RwDg5tffBTbeO8WJ3XHoybNomx/v+8fjxh/jmSeUByPHoI8xiPLGPNh7EN40uAM680Qou9bTwfv8
6HwjbiF4QXCoNyz/Z+pUCm8Hp3rGtgP7AQFreHcu9sLLUS49w5ElcBHofTeUr1BwRExvJCqWjpH5
WD7Q8vZ+1WA08DVH4s8K9zXJXCHNqcZoCEOxHDm7AlYFJeZ34DwH4LLIFL8hZk/Q4sCvi2I4hfHG
TWEPig52KUswzG/GeQj3CnO24BhuXoNyWc3sKJ8iCa1ZTQUrkHMMedErWCnbXCsK+E2rVE6gpzFG
jlleq6TtR/eIfkl8R65caXsloYlmItY5FUb9r7u1MgC+9Ddhrqz/KXwybYOITdOKurhP4Ua/rmcY
ZMwaDNj1GPkPqTAxQf+SdEgfJaZDNBhLRrAIRqujLbGHfa3wgUJf8RDh1sI1n4u4xPxjBpBQcQ58
CvzPAgPk7Jo7znrVU+N/K3B1utJ9LGuKLIDj8EmlDWJ+3t/5e8qU7z6Gif3++/5CETqELs+zqXqF
amFunkYcUkrBwJ9JadUge+zmJEYI/FIaRIUao8McdcZROqX2CLXgz4YSKvBvMgCm2vCosVMdRVH+
qd+SilLLsRBndDoAfwoRqT00z96lOLEmtkeUqmxmjr3850SHtpjjygpYf48ciKq4j/4IEx1QZRuu
uMMTXahRCXvV6Nz2PquFIVHkvZIJs92pxDcQH8aOvPv8BLpMxapmnN+1HmJlZqs1xx+6LFw2N/gR
NCirm5Lvzb48mut97rqYt2MI7aeNjvqAl3loaHFaHYGYbq5HPfHYgn+hBCdZYVjE6EopINRrmJ2Z
Pd6DKv3qhUoGoPv8dL5wGv7CN/AwXj8uRENZvef+m/CYNdWrdQ044Y+Tma8r5assZ42iuKdCIAET
2wy+xl5i0G9BknlISXKwVh8hsM7uOz4bWS+9KvtAQXX+6geUIX1xwnzVlY5G9paOJ+iZqxW8HSVz
ALvkkC4MkPq5GLf5KYUZUQGeDIIjXRe2bndR6u6OpAFUAPW2znWkBfph4khFRIPhKhpleupIf1Ek
nuLvnEg0d6xFpEYxMamLsfq8RcafjBRL3CiTLssb9UxM4kie7Jp3s7Ss9JpFXx0zrr78uKkyiSVy
zrYBdbreCl4dHqlz1BOVHklfUgRKle/FgvSIAUIm7pNEyjyu+mVtqrSOdicS8/92teN28072bTq6
L1FTjn5Xrlctj48oJb7r8EaF8Rc5EH69ao9SlOy8Hyo7QyW+ek5AoEBxEb9372a1B5tlz4v4Nv/y
u4tykEhr5TDY6SKMMedVwkrum5HLdwI2oTDKxhPesRQVYFlcgUTItofvZKc0GYoSnhLqHV5Dp7EI
prlXoV9MJHQo8aLtYDpI0wNcRYow5COYG2toMXZwqZ/9KGY2rj0p3/k/1FvlIb3ur7Q7yiwMVnCt
O0ITCniGtqA4ZY4Ox3ilYFiJ0d2cCuBQdjT+2rqS+S2JgJq3hWSqtDNFL1aKy3vX7oOekMCrV11k
9k2rzn3HOkPULqj9N+B7hgG+TcRN+QMq7aFgy5lcFCZsbK0lhsgGOdxLGDs4pjijr0/tqz76pO+K
YuBDwkx2zeY+LWZI6/mQlm3S8dTvAw48n0MiqGX4sOeAmDXtJFgSI/jMXAFjWGKIVs5of9sSaVWc
OZjWGIdbOV2PMPkf76p8o14X9sdtfjOIaY9zt1suDdADUUyev77mpue7VGc7nuUeL54AwxMWD5Df
rJgeaimNpMXJ50RA3mXTCJKukit3baWJhw+NkWi2i+joBdgI2TZRndtzDs54t3ZNcHsLr6xXooAT
HtQqPr8EZsJJ6Yt2qqu0XIXYHVv5C2yYTqwwZgFUUFf45KrDV9rl2D9+K8qdBljeDmJqZsuqfvkD
hA43nNE+iMvKJ7xp32Rf6Koei5JF4EGlVgAZ/o82AN5BCtKuHycNPZyN8Ff4hkUGqFojn4OdtDN7
lOvQrU3qsn+78b6wC+MThH65/qzzpmf32KwXMquvt7VPwzIjt/nop7AoWaTjbRpv43k4UJ6aeg7J
p6sX06QxQeN3K4kwy4nU0PCHARK2iU04OyCcUJZpMV3nQ2W/YfXEYf2EHZqoMCHeblWmy0oSfx5H
ow2HhmkuD7xapDIHccs6OZ+vwuyvILX7ipOKPXqxYWAbYPpYZgzrNptnGY5D/fJgGIfmXk2lLKG0
OfX+CpGMDPq5gdx0SQwb9PWsJpx2HN7SkJ7KVWMck+KEBlLD4kDhPj2uTNMMjQQwADIjSU3qau4L
BlMXs8tAR4TjIfxSBr9QsztLQ0whLYss+ORSO1LUAwnxt4TjVS2luhmStLp9qCsFQLewIikuV6YT
yEnzi1bsBabmsK+wc7jSHLEyV5SjyyhDkBTrt5HWSk9YETJTZUNW2JxL2EoOFYbeImr5kdBuI3Lx
5PKiyQizzkHuSkx526KoSYAcwTFH2fq33h5WPQBUZzMZFTc7pyDbF2P+Jqigkirz+NcpppAknhzq
1iSKAYFqd67im2V4gK9KOgMmCWo6rJLMA8ZaDqPY55ilAOP+ql7LLSAz6IdfaLNPFy20SBK1RM01
fv2pTSnkWUTJPXWh4Q4JOEK/Qn+9C48Mgn3HwFxYqoH/3D1ecXTDu/+v/d+t6ElsCvfySuu6/Rpm
t5fZgIoTUuHBRbrFe+EEze4oF5s0Y+4oabX2sMlveqzD3prtE9xIrrURv6UZKI2GkDeqnUKBmhK7
JWcCsMDuggZK4DcnQ8jTOR0ZbR6gNexFsaURQ/K1f7+FMyS/dPj2O2EZjkeT80Jp2JjvumMeo7LE
vL5wUEB+5WTjUPGh23rugw2zr4/bEEwntg4nAe5k1Cdc7eHC7My+Dq+bZ78k1LwjcCJov6oyRmVw
rN0NL9ymEQRI3Nc7QP7ySaR99He0UPrOJKtlaEoYiIxrRLg5DzNCiL0QjVJ5myTza8+ZP7Pj5B6Q
p1G5bqTjzjz7jIw8I26NQLVZNDSTji4gJC9UbscFuiORKMwhW8PpIyFt06BEhjIAnfdGZ3hzRNMj
Xm4byRmjjtfJheadTa73WxkpPHeJeFaoXuCkd4yykpdJ2sEjRspSA9tIilZTuWRZ/qaW034nUFRY
8vp/2r2RsCHZksmISBk50RiKTR5ke5g68LbLwgBXimtD+vDDN5+UVg20N8pPQFhl5htEgw11ZKrI
vwiADU7jwIhpRqUY/RBMd3va06+XLyuv4krlROFquh2VTlo+JIEDdYQH9Itx9NFzNtGwND1LQ6UY
9I+K8yp/boAQJIXXOlTv8xQei9WoSabNh1tME6gWaf1fGP22Q89FAz9wUs0f5TNxXZk6kXvvOmKX
/sIKKpif5roNOcW4GymiQaRw18drcC4dH0PzctTICwZevUgXafDQh8D2Ei355oIx8n1+cUy5mXyN
gmE1Q5cFqdoE/xfRUra6218TZaTWgILqpB7bKQnEkPweabB+KUp0iRLLNUTPKKopqjvufmHVtKhO
LSCCkRwPgr6wuxnxxReGcBn+yZMB8qCes+6fVPnjSpZEDzWvw490L7JqtLyNkkcM5VJagaVJvhcm
x6srRcM9+wERg1XpKlZejS0rPbe8u62Q/GYZO15DxSsLqzdItd7SrFXPC5Gwzvv8+cyjAWfB/wyb
5sMXlOBHIYNwRcvM/lXMvwAkK9pJ4A79+OCUhiF3CGXv6meUgNyOeFZESqOSpWB/3UsP9x5H+EKp
rcFlydzYBnce0zUj1YlP1HLDTwKVCQWRDRE8sjDhu7PYA66f8kAZsj8S/8TqWi/DGOwiPiSmmR5t
rn3401auHg/Uekht6JpwC8unRADUbQSiO0DR+nx4sGL9sc7M26dHZOeqWmZIvxvsohOytJSugfNb
RqUL3792frO43lgTabWkUC4xsbod6lvXbpoDi0ApdF7O9+e6FMiAOJUtgmQ7oEf6XmN8G5PYIcN0
TOUJhVqAJmNwhBvSS+xDeUfwGyVBbQ1fj4HolCnhXrZ5UCxpA+7/hrSM4sikX3rPtqr1RhfNlcuY
YD4IGApNyBSPCqaqtfFH7LZ7q6sBSyaJD7wgSDAUO3j0TQ5cHkh24fp3a1ufm/MP8Hocw4xdFPw5
yom7fymAeLJ0pPhVq3IjWAdXcrNqY+BcKJTO8nKcnH4N6HLoMo4sXyRmy5KwioiYl5a6uYipBb4F
TCyQ/nx/I8cMHk2A0LMGhqHPL9NoHiyv5LKqWBmLP/Qjcnp4+KqZvAZvGGyz40p3R+ca51/6lF94
1Wn8xA6oj/IdXvV2rag4gdH4wgZEMl8bgPBMJoEqJSufGUntAfBWRJL7FLvhLNPBa+nz3MZtvSau
LBfiZKy1V7XPPq0KFNZErDgO6o83wo9x58SCfkuDDI28J6+Cu6HKjjqmq1Our/qHWMeQjKDGMziE
4BXHgjlQXd7IXxIPzf4ynfWpN2GyaLFQkTSlrjR06pA/jFY4whj+7l5Jgi0vt2BCDuRbk1ePhSPw
m3hwJp77sOrRVtIks9t+uxe3z7CmdrbaLYufykqNFaNx57WlGuj8sdX4jhT7MD5JHygG6TVdQQjb
1rDfMC20ZhSdMZ94Gi6stsmDSI6pS6MR7cunaBUgzwqrWC8Q/wulo6SEUi0scdmt/v+VlpXDWCHi
0RZDTDNDBZQYrrxsrk6CRX4fNoOqVMssKynm/HTHy1zxi0K6I1c8+mDbzHfgHkNfOu2IUk/3DICo
mPvOMAlolTLfZwPBJhJMcDshIUijvipZ8maxT86r36wSrDMQFodtMoz+GQmlyHf/TaD6Nv2lnx8J
Roj9CAIO8bb9KqJ6PquFvBWljAhTEw9agmWQMvpmCp2G/j17g0ttWPO4QG6IKmIfvkhI3q3ZAGwS
GlYVqwLymwM3+g2eQJHs/++RF4AD24sXbWi1g1VTpUDi1qbINixYGhvJ+ahQjejVDeqL2wvMfaQ2
313kqNq+bxzoaddzum7yPuOTCAoMA/wiXnSLc8QPFLQVvzOehNyghkR8x60HPzHWZTqmlTbturBw
wR77E4qcAj656H5Ey4my3wxgz2uxfdH6n+YIMpgMipaa16vG1InpPYYBku7xNiczjxc1EQ7LIYdd
GJ+xlqFG2JQoxdJmLrAJ1cGZpLxaD295gWgTjqj9rDB4OVwMyyKhCXxECW6x0QxPGmVvB5qVOwzd
9Mjlv8w4PmOQAXrkJ7KEdEAwmm8ZnUReb/HLkrvnQwrXSl9wY9HMV7DYmo4EbNE5tdR34+pikGwR
11W7hsGW50EPoGJyfytqGYqVvtD3QBNSqc9bJbQYDMQ1p7LX4e/02nBEfj+kYYIMIbgcEDVCG2C4
KhceSqeQ61ZMTbOYkvtVRkcQZ97jVfJZatOhkqyVvs+RJp3pD1NNFXpP3xpV9r/SzgAUIsetXMBg
m39BveONEregkI02p9tGIgKe8u3pOewdMaHE4FA0XABiIAlFJ/5LgqZrcH7O0FsHbLx/gIqyRU2G
oPo+cg/HTOhHBs913rGjWasKfFU+jibbAk3OFKK0+SBZ+a2lxc6DxE4EiNi7yUS20epw9jyc4PKt
LpsIJi5cdWpk9k6p6R1N4Myb5cgL24Unzv8mPCSsqkALNFrVBFvalejkXM1Q9PnPCgt1NWDAczlZ
D2JZA9PMvDj0HCYe5eDPGyLZTOO9rMMtJrnVcPllxySDNy61siO2TY2D7U8/rgfJZPdC5h8isfHe
yyxp1IAzKS6CImIuez1dM18T7J58TjF/kBXfCsk462hKu9NjxI61xiDCn241SuG9/vBAsbzB3B/y
Hrq/Afzd/7M7vFQbwIasrzW0TUUHY2vt6V3s5sr/3NgmAD+ANspMl/ylIX1eIBgpVTbLNH8FYiZg
bEqsv/bp2ZF85eVZZQ5XJayP9Cwc++IFzAjhW9P/OREeoOYEWlbv9ZuhtzNWaMs5PHxIqyaHwR8K
qmR7HdCoFpGbhQ7ZfYaPzzDTNqlIbCmYlkcpAWpE6wdqhb+BEE/3vryNCbKsn8dIqUpAu/vg0yjA
paOG4JzC2jG/4RvjwkFRSuan+qL2gk9Vibi4uDkyjS4ER8XaysqoC8XBqbKWbwquUop6dO9czmfw
vfkm/Fec4J63KNEyzKUDtJHawGnUN9PUtjGiqF9lLWY0IU9yOu+R3oQO3B0vHj8QLcK3qNOWJgb1
dOWGIrIfb7ZCqphPFxI2VtubxaTe3INepf8lwKvDkivxxkOxnIFovUcpV5SThEUR3xkeqcpyI3A/
+AFhj1n7xan00y0q2XZAKiEeOusNtSXxD3m68fVRwEhnjoYT7/k7kjLJpHK5F03R1cJpZ9aQHDbC
gCMfA9RnnBb3zMm3LNc52hykWzTz2OLKU7JgarES+ZEN6eHTyPoKMP2f0CndmBERmZF+wW3ri48V
hHw906ZnM58f74tJBBPqKGF1oX9qaqVul8S91aCyQgcPj2t9Ta3VrNC9GUZk9QBCEZRKEqd0iR0R
sgYIOwpY++yZhXX8H9W6QQSfDNe4jFk9QEvEHUdNxBL0LhQ8NT4+9BaeydziV018oBr6RdgjQ3HZ
xnGU76XsWnLy8XSW1SGBzSCq8A8Wo8Vg5SPYsUjdKA9An1N/X6I0r8EgYyaOcDxnqx78FOGxlMYi
/2m13N1BHRVLkjwzpjIiudAoZ6O6e2LWEY5K0V9lispogqGZq77gyKOd5nr4cmgcngCR01fXMc6G
1G3jp82cwJv2LyDcGRhSMKrvim/PuYvG3sXA09Jhcxo9rDAXzkaWasshZAEevdKTJsQigqxhqhso
1ZLXguepwxgqdif9u0gCFVE4A2JcYNA1NVo39eDmFKolnHE8N/yN38ilv5vXfzA2QDD5NVrk+jxb
sxBI5YBMha3qeXvr4fnFHFg9uAq12HdfLT7877+pJ0xIiMdCuFyP398DJIM8BUHiG5G9Omr4Ju6f
0y83lZ8Z/Qw1HpLTdj6ML79NhKZcmAildABA8hmvMQiKSgClykGq+zYQdkYZAE0nNENtQoJZ8KDB
hPkQLtOQ1b8G9rGgSHfZC1cDD+iUTT5Bvrj5xfyg7MLtyoIPIBqpFURtEYG10tAZqFI76V9HqKqX
1nP6oBMpGsL3g01YT5+s6Y2k8KxlMdOBUI94eLalNGTYEsW95uYHA9xMJrevJPr6WPCeJUmHGUWh
r4lgDvJQZuwcS7X4VShQ4RDwotgLSOYiPPmZi6Ebi11fs0tmG5mcZ0+Qa213ayrEynEemA4tJLd/
XoQfe22UuzIUNpB6WwXDWGtKyPIQ4O6KXJkNBtca35MoBOppSSr3yEtmr0iGCKF+S7NeuNMhjTkV
rl7s9XW19FP++TFg5cHIQtS38QJ3KNionZi1gYj1VPBNhCW5Nv5qLLvd+l9a2SHEGkscQNl+zk/4
BHsylLFn7LjrHw7L0QM3/c4hVxS7fMARPYKAiRIJp6k9a8/BOhTYWkPeLaCkJK76LlF1G8fz77WL
Vih3uOh0ZwyvsnDN0e18XyCPnT3vNpZ8ceUrLRSS0RP+gBUnKB172th9sw/lpRt6+kFtPuqq9wTZ
DurN2XEPOlVbWO/vYayfrSfQTWkGAvhQBCO6rkMgpXYl7W4r4P6Kip2CAvNIR6Ngq3TnOVZlsB3b
XppDej5yfirfvymICrvlesu1lyMPZqalMNO1dkNC0D43IhsE560rIWW995aftDeOh8olin32G48Z
PKTTDuEm9ScFbK+OMxX4jrqTkb652zTJog2nIlgnVjR48ytuVuFLdH1/DiiZaeAzJwMY3asllDV5
vhDncDumBP9WU/LvrHGKgas5Roe5kO9a2F1CkHFyGrELg3wAQ+H5AUysYXndaVVG9/eFsJgdqgtf
6tJEBy6/7/uS9XexujH8hkTcp0w/sIAzr2E5OzzPZ5pA6ZxQhs/Upl3/rQIyvQTot1/W5n2MXwiy
UBxAuWjgnoFy/7NgS2z8rQ8XoUC8RTUmxfeoaIGsrhiOXU3QbRcJWUZQFn61MNOlp5wec7xL1M1d
XYb/e5jqH4iIwk3qytaUl6BJB0OEbDCJhw3xl0+GEuAZ9ER4nEEHmNQ5S6i0Y2rik+vv633LU29P
QqMGpzxfKlu7wrT1NPs4q0Rwk1Bbj1Bwxr7xwuUyukwk+d2/yi0xD8OwPbHonATdj9SSGMuaS1k+
2ZPaP7DYu2lE36AZGZMTUy/GlDJ5nYOxCHyzpTIlAOdDqW+a954+POxPlE63+8VBY3o7GV8xBRwG
pNcnGafPjqxkOFUIbqLC71VAvRasHqjspNsiWP9yQ3r9tYiX0/MqisE2o3ub0/CSQSswZm2FiU40
wj3VV5PeePAjuc9keiCRt5ETn3/x5sDD0pWRF8+eefR9TJu6aEiEJQC5TDJugq4vcBHaNOCzo/tJ
ujlQZLj47d052QwdgvZDurOM2sz3FcQ36uZ1jMTiQImG45Yo2dwsgfjy3wNUwL6XpDLuWviUo3vB
39O1DvduatmwpIEAQkE1rN+Sth3zPcjJJ2yAMSisktljDwrPYWdGLSjdzjIihaMia6Dk+oP9XhBi
6TCdJB9yq/HQQ8K96b94/sxGACPR71+clmeDUx8OB+hUT5FQuG6S+9S1boCl5m11P0mvcO3z2ROD
iiVLUjyGAQ+cmmno60Xw+LK4CimGIVzv2jdHBzirhrS53R9tdfpUJd04/TVN//Bv6dVTEgVdc+xr
5xONi9BkSvliOxNM2n0biGIVCN68zhZZH/Ndg7FOcTjNUGoN/y0BwCQm1NIyyN8eN8HKM7dGfNMr
0SEPNCIfc45yzI8YDxsmy9oyfK5DfTE/IYb8mszy6WCqkJZ5QAvbaFvt5In4+SkRz0ehElUy+eUZ
LwWyqch8PrlwwCK89dG7N0YRZ1ub14II+9uG3jbAVT88YORG6VN4lUdgM3tAbIfBNvbcntYfAD6r
XI9zCZX/qI2w3NhvvnBDJmfZqv99eFVM+5QiC1s1iLjL43HTYqcrwgxZkVpm8xXdb4of2nMWu+iQ
npFs0shEglYonGhQ9CX236yqTq8yzvjAWzOc4SVnk/MeDazPh+XrAF09oc8o8eKRGmwS8AEOwlCZ
IseSROwgAOckJc0kmOcTW4bIaY4lUfgYNerROqT5QjO9xKE0jAHipZJ6EYKwBxzVJWOczsZTCAKG
QUHEJTUgA72uB8F0NlU5RjHs9q96tV8Z6DvwU6Aw1f986Vl+lQ958QFGAxFI/VgURImUw4fTLBZ5
46l8DzzWG+Byn4Ml0hAXjn/zt3m3fc/A1idfvS9EK8p8Vw+l/2bQEiLapFV4kPueNKXnofZZaazM
O3M6PChz7e6aso/EgFUrOGLPINTjLs5BGKDLb1yBAajPwJnyaw3mfFFS2pSMwVYOXDhywZGCrI+J
dmKqtHF23LdmTsvrVjaS/cR/VwP7ezARpZW7xgBVMMnS/Lc6FhWitume1Mmg/IeXC32nVlozU2tw
ZpFuE5nNf3B9PhnimJKHmnAH2kP8HuRt6F5WPvYGITBeMFMggKNS/CCiZspPaUV3/XE/gbYeHPmW
c3SDJpFsDtW6fa2ws7J5VHPTqBwpXySBWeTp30l1+SV2yP3WXrscZKxTAAaXghmLLQzieOT/qt/R
6OsDpkxUDfxq6Gmc0aNXosMXifiOHHfznM+W5RqrUKSV32Q66hvoQz9fbKFhVodUl8/f72YR507o
ktoYuz/vPuzA883w+6dLVmx2bzcUTzziNsJcVnTKvELS3vFIUUW1YZrFSqanW0p/3EwG6cMf4goC
bFtTr6nvidlS23sB+TO8wO7Bt0KVgae/asH4VO6LVg3Rqy6ZqyOZiEGYTYdP1gvHzE/WItyvgoD5
uthMVvTUd+0kSggnDxSB3I94Adp4WHAGztj7lzRucD67EdKb8+bu6Sz+Y8CouA8Fd5cVgpw4TXj4
dW7Dai5r1cEuiDuj35iX4LE57JTPbsdXCuHDB3WBQotZfc8mda929fycVRKuhgqnLOoTZwxfEFJm
IKua9EyccUU8QOn5m+yiydr+UEI/nFA70l3431kV0X0Hc6OyY71dobdNt2dtxq3rhPQukS3yNshu
WWmSpzj31tjZRJO1FFY/Z+yDwJ0umbO6udCdpmCNjjH3hs3OvpGR4tZuuz66Et0DQvQSlpjT8UtS
tSvBU+Jphw8dfxNcZzP137CveeyDJefrgUsy8jkaeGrmCJBUmUdonm6ip6F+6dm4DLEa1BYBVAlO
ePFCM2cnAkP5ViNhnThXYOwHq9Wah629vC4rau4KhCHwSpmiD/JjBLz6GrpKF+jwts27hISDAtga
gq+HGR9EWby1QDAXqOLGul2uJ4NeP3Z0b9QSLVlFy/GP20SXDHmVk5e7de9HIt+jhv1Qpq2cdxtg
E3MXR/ZE1up48M4np9OIXb4eTR63vgV2gvlySZR8KjqvCQjs60BG/433UBDoJc5JBI2z3Jwsb2fz
RD2ThasxgvreOVwF/ULf6Wg2nS8uNhPJqYru96WbNn+5YxZcbkvRXf5aqARBnfNBQY83MG7Njhy2
/GGZbJS4eoKi+9neyl7jWdeFUcnkKsGkhMByw999TNGCtzk7HcdsUz13/2dGLChVvNw0yZtdKRg2
P36tv8jBHhxS5s+KdndB6ifQ+lw8+Ix1aVgOyKq6FyTqb/RstjumH24yMcf7sg1PoCBdsTyC4CMl
UTr4Cjs/Ej51z3+4kFm/plVzLZC71MCx8jVAxH0sX8ASASyiPiS4KlOU3DvFLcSQdkv4kwXd+TQq
xYzEbGY71sVc9hmwsGqzF+X65mETj/iH/oii2o/EakoayB2SzabOXE/2JqtAX/uLDSxrR/vbri+l
9f1YDktoq1ohXwMzJbEqWoGqZrBnGOOWoLqVB8KXVU+vHdjz16ZrvmKud2hLe3ZvQuvytupQEpzM
orbVWiakfi5ftda2fMTrsnKZ7YyoPGlmp8a0ThjdyQEHQWwZv9ukoV++lW9BejtrLKTx/xdN4hIU
tOY5b1N03rzqmsI55++fH/+I/YMW2utkmn/OlrkNiLcfvKVKY8eUjeJPUdHRtKnXwda97wEDQ8pF
qacSBpMqMLIB+JaZHRhXko+rZXLOhreJHxePlatDIjPAxqCREzQSsjcfLmg6EfZv5y4koSC+zZZ5
bgZ4PPozGBSk0A8ykf//VZVUqaoUwuqd4EH5OwYQR4f0cFRbjfxcA9lB2PU8FVfP+1yNGefqdDNH
F2hn01b2c4OlOWw575Iqa7B6w/UzXHs6ltbv13NjS3dYxzOYYtoLjJTWzyMZI/LfLbdFQ+Kj9a1g
sDiNLb5WbDF7I1b/oT3o+qvRF/X5E0rKFwP48c8uWes0jki9kEv0xwau2hVM0htEEsJbCx9b++1Y
uTrIA5aPa+6uMVkdYQuTjoRtkpq4qauJpXDAMjWkT70TAbKXanzbkTols9M/NfhoNbKPpNbnedwL
cSeQ/q5nUvzPmU2djve5b9atiUJWGnLToLE8nrvfwFSY10vPeJTj0uNx9OoGLyLDe2vV+NG6eAVm
/cMbvmmc/2AerOCJ5lMLmwuh60MDLepL/nTMcEu1LKmRCYMrgupc9xskTz69orYFEdm2jUr/Iah4
H2y8oY7DkDDAsmND8oQxzHxgF7zd0J4HVEcEAjoNOTpK64AGKZfAvsN4KFBRR/REPXJFqweKQXYR
2OiDVzVyLoWql/R9cczPT+Kqi/ksLXUh2ePpw3UVXmKpBllShFviFHyWRl9jllsZYTHHPHO35Anf
ata0L7UnQ1kH7uTjptZ2lANJ3OwgZNzKtdHlPKsYD976EKAEsnSMLcrSIikceul4VvbWDOUx2hBD
cPXrb8m/R3rGQa3XhLTcjBqB543DZhzq1vdGnOoYNWBKUwx6AhtETtQorP3RY5AVRtNnpvRFpFLo
GlJp6ukWysb6dnlucGcUWyBIfRjwfTMCXbVnhEzzwQNOFHQAE+MwIsGVdMBCPN4pZL0CZuMUGGPp
8M3OHIs7lu8qYc2pOcHzmo3d0TAfcIk7uacm7dyeVZ+lL7DVJ5J7rt3yZmme3amThA7nRu7nGoQA
pPE2DWlY+lizgIm9hRFG3lqlUrGTR4Wluf3zA1JkINhM3pq7oqHJSDlNsFJT6PAb9B1RQ/utkYe/
VDy1RUhjEAg1seuxDyG08y/1weVpZnJuzl4iHzUzuTLlCRfIMAbktppVElIq9aJBX9Zs+GxU+EIY
G2bfeStAkRgQ8+SCsQuNmBMSF2o/CAQmqtRKAmqfpE0PMQDeh2dpFrf/pXFnPpCVbAX9SKwPL5Qe
ZAtzDMWvl4fwH2LJN/NEWFnp29DHhP+f4ifACScGMb5BRo7wRQkZhKDo8MVkAe4mTbTcdRBdvLJB
+2CB7I6AL4IJ8RFG6YXhJzTlmMts7eu0t29h7mxFOA2PTrDJtRm9pKT3XE3gPmCowVawWdHOQcEQ
EwdI1W6uRZlcsaJvlmu2FHtE1nNAnCLIlKqV9OFcyEnaC63g8VLF236aSAROdST62Ngwd/iACond
vZAJgLJMrAi6vVimxZ51na71sej8ueC+USem1c/2MLnMf669oGmIfzP55XWwzs8qOvpc5Seumz/k
WM48z3DzHcD5LrQYKJPcub+vHzg5cvunjrf2hb9aSIdAwlM2RAyHt4OS6YK4eJa5AlOpzGHo5qhA
1eS44KAeNk/EaYbJ6el/G/s+QVU7+G7RaJQ2Z6GV7eziIGWF7wJVXRQuiCbJk3MpprKuUek258fF
znTyxEYsN2cZFx86Xlu8Fh7LogtZYEKHEzdEFFtd8ehChDtbDheyMhf3gLodLuibDjsP3TVur1BB
wmEfpaJSob9LjbUKFpk+4VthWt2xmyqxhrh64z03D/MRzMtOOI9P9Yh3IUi367cY9fPTbWjJ6Vvg
bcph47vV+ZApvqPd0nwI5jRzV8BYUIMu/RFVnjiIw88uINlxn2aH3xfWhQlArrcYMete0dYXZ0E3
Jh7rmZP07A9BSFiwhcdAWbtxT9CB1oxkQTdUB2/4ArZFUD4hDN71pGh0hrjS+iQGVWgDTE+cmf01
F/9Jg7eDY/vpV1P7q3edUNt52iqCa24UysNaEF74UM0sf05xiVkihI0x+MoOjMyHuTuqeAbSLDY9
l/tVNRYpHoDoRGusyo8tcuhu+UpX1tB0wwacelOdajvbu0MYEBeD1AHwtl4rh9ozdSj8l7cAgDyk
TVfIVomvMD93JIYWXnzdLL2CNhYp7QIOv6UsIVCBZCHyJGLJ5UqTiAblzLp1u68UGArDbqRfQb8N
LEn3cvS3CZOHBBSjgK7+v1VkcJUQuashQMbvMFKpbeqok30etwTaofgmCsvPmN0Pkv7bpqc7cYqY
EOkX7doy44Sgl2TPcjq+4CvNjavj2iAf4jqEk07OVPGPqCbWd6HwXl8tqiPCsStg804G7VFaUZ9j
aCyEP3H7w8NRId9aqH8GXHVWVTFdXkjuiiSfrCC2zzO/hiUGp7R1Ut9lWsmLYGtk8ueOfw3m2aur
EWL8x5013ZWj5ZGOVfYWZGqMMYcjHOYAfnXOH9yQhyCYdxy/MD7UV1tn8j4HcGb9a95IHeE7uiQm
0jw+8tgSsEwy0h9pQaYfhN2R4Mj07pyC+c3YbBgEbf5ImFo8pLgZNue5gJBZNcPW2CwHPYcLHTqv
pWGjl4tQWcbj9l3hPRc23J1ieq2VSQ/3z2jEyNTyEzMmOhHF5tSe9rs6no67CKH9xwSYGxroYXQQ
GVye0fWcI6XbUSajGSYSSOfD6NeK1hFdUFouZZFhVjLvH9NwdJ9i53wsbCG0cpE1vT/mwtf1kKGN
ZONc3GB/T4fZpaZKOshEOUPkvBUQ/xPEpVrBAzyzn8DhxxOvVkqU2qaCtUlPPold8gRflSicFhTf
k6m4p6EKHVxD51/BNI+FK6ibpJdvTcjbO9/EBgrh5DRSwAqBe1HFJBz5XC9xDwEc7WgQ+w+nO9jI
BTa87MXOYclpi1PTrQbtAuO75TagQPuGk6LFO6FZMOculw4O1KJWo6N8+w488wZ9RrGteUsTSCF8
dV1tu0jLvlDpFyUJS6oXgzVUtMRmk1Iz03zvRcIw/iKgNdONUp/ss7TBDpwQGHcaKu5lj4uodTbD
RsahI8QU3ykKo3hjiuA8LfnPgdL3ViLrJbIvy0dDKpJQ1VFaO5HI3z78jkhIvjimqk6ga+HEJbnN
jDu5Xa/ml3Z3A6xyUIcd1Khfd5ZEZgFvl0PN7TU3ePriEMc7vcw005AynrD0qfe8t02a8XXApvb/
Dm4+uvGdM1RNl2JMETuhWwu4o1mp0UYCSb/0LRX1tj+p98kgjx0POwODdtEYwSA2nI5cuEvIUSGI
nsWMMObh56MJ/QhzRq8mbjrAsUP7oD3kqznPDu9vb3E9sMddP7LCCA5kjSyR3Zp7rJmAgR5jwNUf
pHb6h6Jpxyneiyepw97r3wnbvQ8Ag4XncNRrN95uxmTodtMjg8SLz8qdW/ViFTZOVRVnHz1yJh7l
lh3MYUXyDR6P5LPma2Q+h0sE8XFXMxzES8fW5tug2nWWtrHC6h6PppOaMYxs4bp6zhv/dq9FLmE0
vH4RaarH6/0aD08qyg3E8zcY0Nc3te5IbBEhW+CsfwE7N7fJ2NOIU0LuS+DmM7SNVFFuGYqjqIYp
hz5TJ8C/DyvgM7CYp/a8hjr4qIfOR5ZzLES1Vb0u1WNuNWoZ6OsvJ2Sg0jfAbBvlGcMmLfX9tRtg
HcMvKzMV1ZgRIylHd8V23MV1P36JebJGjnZIGzgkdbCsnkDi2UvYKc6OZyGqflVVyggSz/9lhPUl
HeAphBhc2GPrq12cIlXAYDJttt7TOo1PPtseDegFNahwsYUYFh8WC0HvMnc+nzALEL5Bp0/l4E4B
5kdQ1ImKfF7bCUX71w4X/8rqNuC9t4humkSewAe7sU5zL+oKNTsw4+j2Xm+1Lpg5nwKfjAoR0ijx
CCdCmSVaPQf1N9zFWSNXXZ/gblwDOj6ff8PhdOjAWA00AYxHnkos0tx9PA4L8Llcv/onCmp+a+kr
KXdFlGNt36tFNTKuSDi3qfJo8F71FDQHRO9hrGXCCii+smvCfb64+8PA5g4pX/v3c6KxQ40Xb6xv
Pv7c0X02m0Jw9Tr8oeAjjQNx3oRpEYi7Jfe3Z6XRPs4S2G/Ol41+8RyHwcy7COBd4KkwvtKiCHVL
v91cPuHFR+2BxP/uqB0iS2GNccgGTLtoE2kBU2djeos+ibadFqBRnEfBqD7SJajrxPRRLhHcP49M
mPBDIoBdkw6yLvpi0NYT84RsYmRnBoy3dxWmYsxsMDpwsXipjzIOEusTwuBMv3WL6PaOy/GuUH4J
4lQNl1alN3Yh0i0l4l1hXA5KG6NLVJXr2XCv5rlJEM5DJN8/UKZgQo2yKZSaRDwqT2z2rVug6n6A
5eqKUoOjvxS7i04gvR8X7MQ6OXOXXb2mul3EsOOSHcNXs7QhZVHYIYnpmnFfXUikSdOrk2CWpaUO
GgKLIPN6tCMrBm34AfysWBM7pURezmltRfsw+7r5NkjrDjHgtPjq2t4tW/oBFj1lGYe9QLdTEmEn
9TDLwJvb2h4jtU57rXYL5gbd6caDF76ZYEEgDQJNszBC3ihlr77zferILJwFqHOmpQ3Zx/pkA47U
ifmb3FyR1qxNJPg+eN2YXZF4E/bCwuiCZqDIdNWESp/q150p25Kg/3/DaEmJQcBVjoTg68O+/9CS
MctU3YIfoArCn7FzsOv+wY6y885ZGCTD0VrPXl8ehuqarA6Nb5AkEKpcgKDrAZPgXsrvKEdCqOeB
CKDjmnjomFc/EPo3u4S49Iz5dHZoZ8dH4XKVmjnIfjxJO3xIunpLFvCclSEOEn+rm7NJIWoFbuIh
FX+DOWg/Hljv0nXT6NFwVTzDFaqpYmv9apjh22cT7v8KBa9wbNIl0Qnamso64qG1ZU0paGrt8aAD
yzjzs8/QHq0W6vUPvDp2V/d2nSE7VsDdKxSdkmJVJPXYn8z8SsVbhb6BC9cDKrNbFFnSGZy26btp
ks2FpoOBO0AurTc9hCfoA97sJ7AA/0KjFHJFyWkDSs87dFqMEwcbYHcPFMEUKdeVTB+7/55dFQkf
2I9cg8DLIwf86IEQszgzCM4BeCI5mB/+3g91O2vO+NnkTKoZOGWyz5XnCKhvFvL3CueG44Iys2tj
kSRmmZIrHA0/703FIxD5p+66M40k43sgM54l9jSAUiD4wtsx503JSCP66qjp9lTux5IYcHliLuOn
hS6SgpRnzWg7svJWpca6QXXFCcZuAXNNZUF676WldfMykjO/m0ersAQuoTQhUPjjFQcn1KH7XGi/
L0twtaECpAlNtJs1KJAHPtLMUDF4BWihUobZuOaeXBEpfsSB06dgt1ZucXTrRnGHBnL1M3dT9KfW
g5lKwaQgip181xd5NoSyIOH//c4ypbwx1EWc6PWhvoGOaucGCckXYn2bK5tyrjF4rV4+OPNcWXYG
L3Igc/hwGkpMquXDSl8mQJSBroHGuK0evyRSzmc1+rRbIPi6APygEBejm38HLQelFHrmmFuzVp9s
1AyxDwpoMyVOhm7LBFdFX9/1WlD1YexT+Mqql/9jKkpXq88Qyt/npltF/ISLwER66DsLgpsTNgfj
LAHYA6X/KwZsBfb+YlKiA/QMBEWgLFNY0vUFnx+/ETTDHpFsIt8HOJbh/XlKJbiaDZVCkRYCkook
Kg7rdZh0ylrgnoJVcbUCm7k7tPEijx0R47bt9REu2fyyyaMm8zSJH9nkMGwbuc6ndibp05CAHv0f
AfwF7y3G2XFjA88lu1J3aszwAj56e+bPsN+afEbP5t9MUjVg03kjYTe1sVetJvnkcio4s/YFbMof
fOYRXhslATDIyEJcGHrgvjUS8pjiZh4pQtsE1v8FJYbU9cDH+wI5GdJyV8MnuxxAUiBwPBxYbS+B
t348k3m/7KAgyxaupG9oeiZ6JKA3z7o0Mmu5SrBjmcqbnElSv1HC47bMN5ItnZ/Tokov8mV0A7YE
UOqP19er0N8mFqy8YPnA84I+VjC+lFUtVz0Y5Pv9W1+bdltN4QlLKWF45Q9qqeDR0bhJw7Nzel6o
FoAxWIPAp+Wl7uH+V64Rl/s0m2fvgo28FeKhX6KOuk4MpMYuS8s6oviXHy2WOeS7TLb4BAgQimKU
5jxjhlVaZBOEWgGzufHrwvBBBDoSm5xZc/XpQlE+MTGcVsqvmhDNzea0PT+9K649LKkq2J4X7L08
Mm9dYaq96W54bCB5YHibXWobk5FiExtvSljnyxGxTfpI3rC1NffysBhyQwJSuZf7sUP60nQzVFK3
87jUAwir/TDX4whkaLZuY8ItFuN/Hv0X3Jwj+Nq8TQu+UAdTKuFrwq5xKyycP2lPgvVHqLUjGtBH
1aqNba2YU7zeyKO8crPI1moc9T1wmUCsBtvhtIlkIxcDg0Kt0yPWMt+IGnpjdKmN3F/SNWmJBdEt
CdXzWGjhUIsdTUMFGECO1zjZsPN14J/ghh6HHu1R3XHterZIcLk5w9cRqWTXYzUz8d3H74iGK7Gj
V2PCLr07maAoCiKePaSjPEOjVABvQhDYZbuUDg6/FUyHCQRFNUwDeCen0ycYhRW9nZ6AyEKMOA6E
qFfEaWxpUmIsW5d10a978cg0COM+VqDyfSIzIKULbOy/HZFJ8BFcQxeWeI9aYYpn35TIiO7F4ukP
oKzW2X8teaISfvHCbOG1uiOyzhdvHw5S6zVeFmvZWKXm3252qtX+vUefcqumnxi9/8gcGapkHrMT
MfbVKPxoWIUC1wWRp3AOHzItV8IzOah9dXlXtREX/dIi7bikqi1I3ZNF6reWnTgkJL+RAaMQ/9lj
Zn608drg3WJggzQuV3I0t8KxlJ8wcodF/vfvb/+I5PEw5LOazAsXj1ueNwMJX76tHiwvfKNtShvs
rKFSJyEQXJmRaQYbR3YnxxE8XVLIth/lWbUEvAsthP8LIOtV2Fz2Ra5xuKU8+UAMJ1b4AEiJ1m8n
trLVmhZFCDk9L/u2bmXkAh/8Oefnlw3D/ul1ax2D6QtBUySLPuaDQsJxdXjT4l9FdugGqYpxHWLr
nSWu4UtIBhCJybHp3xM3+n9Pen3ZEgVOURlZPO+cirmkyFo1YChxu6BLC05fHwrCJ5BdYOCD4yF+
sQoDZfMa0M0TkmiPidS7TEE/ULR6JMM7OSRzxVGWzMz4dm3YmXZSU12lPrxqiX0XqXNPcIqUPZRT
AW/j0MBsKnDymBvcHGX8x6poRpiQorOJPQCw4fFzMQ54I5bu1wUj5agXpoE3oRyhIT4utuIYfbrd
wWla87n9shUEdZtsShiWChlOcFLH7FGctQ66sySkWBHnQJlR3Mdbk5QB7E+PU3ooTprOmIK3p1bD
GrtTGWzosb9I59iddk+QUBbnwB77hvvQ73UDJZgORKASM/UiveFfmNC29VBf7tazGVmRbq7r9ZqI
z8hcz8L06+B31hNkAuS9T76QKmovOIyMGb+r3Ym2Qv2ZKGW85215tMX9bV3R5Y7CKA9xgLnjNvID
c8bsqIio/Vut3y4X7NsiObYgNCKbY+LWSMQnCXbDICTk+4w5e5b4ScMG/fWR1OcALAucCLHD2T4h
XUq7g7POmKw1ncOyfOqYbVWWwK6+lrwClZD9EW1J7FE5thJm1nku34Be3b45vFnbzz1bX27P0IVu
rylt2OUj7mmNcMlMAr10Ikl2z+q5CiF4WfHBocdIjc+OGeMKMcuHe0aJ//0m/HGuVS9gDslEic5X
/+bBsj0z7GQfVOHLtUPAGgaRG13vmxhbqK6Y5O7E5qpvs1xwNPQJP6J9TZ/jZz27SMDROL1/6lrR
nuYSfP173qqkRuF6YOZyA7adAGMX4z0Yfd89iSKuZQwcBO3f2GXOHhm91Fk3ZOAKVGlR85lCFLOT
IrN3b8GB4OzilzgK6SX7RLaJsgOlkWmlzVFxZlNrjC0HOIPmE3v+VLBHf13KJ97Zu4tZkzC+4fU/
Il88H5Ih0V9gfr9z//FDMCS9wloNsXb2T8DSUWz1on2whLcnmcuKm01yGvIuXS9DbMe1ZDxI69f7
iYA9I5fhTMqryvsvPB67nJfQ9bW31/tZufMy+TN+N48h7l0LiZqFByz9zw3plH2J4UxIw8jbCcKa
Z5SC11pdz/nU1LvfHydLqF/2CZu41pPT+vPF5314CZQjI/kMFA91bAHBvczEz32FVqR/JwhUUdgS
rDS0oRbRWP/GpJmASrQIHDWOlHJs4+EppjJF9lDRLfK3F1Q5dDjSuN1P4piNPQ6+vbqxkj51A19E
YmYCfgCSX3nPVrVK5h7HyikZ1WEzTp5+zyFK4ZLAXQoAU2Lpk4ODuFkxFZNf/j7b69OJyMAP5M+v
q9ZHHnmUSbDnqjS0FWFV9PC8cVhYGaPcWrjLJRZ4YFgSvDmJKcssvo9oFf8Bty4bdyfcEkk1eC+Z
tmhMHHa+RbNOrpRuM1JUuCzd3S45yyzKziLDruUFwLYZKev3GSkfhQnH64kCefZcCKCclEFwSMd5
b8BqMd0hIAZfNq48BXdX+9zE8pkIe+LKQGET+QeDA8ivXdkxVGxZ9hHds6av3uyUijCotxnh8KY+
TEBHVXZPYk5tVGky/HcclsmcyDjiLmH/nipC2oNZ2/J8JKqzhUmohpuzjTZjj/ajG3tS4hPJre3k
Z1/ONaDFEzZk2cJpeJXShfXaQ1B83yWVCj1ar7zXr4aioKfPrZiX9hFLDxXWTqwxtCQXRyN3iOf9
hdv5eBmSJFQizSdOQm0F6c6AVmmsxVR8wpTEHq5bdFNStHPxoUcAo5vsU+YW/Jdy+iDYDhfb4lPG
FMYk0yxJD5xRrEE5BBFdkRoXGK/GvPWuz9p9qdlDR8GAxss+eXQ8k5XFAYJLJ3TA5pF9LJf40Ika
/8xyW+2ZPcuRKr1c1Y3K5tPaLkQUpRzJ2QEyqCDxDDKDU9YPbuAUGlA0O7hZ6qikhtTffMxtxHh3
X8mTeSoMx7pr2EMtKI2sDsj1uLw7iC4jym83otQaGB1epN5PwhDRATwIkJKYgq+tDUskPm2nIZH7
cP9PjRW2UpXlyvi+xERrb0ru/MysgxMzZ+WJOA8VY63veII431pb+ub0r9yqqLoLU5G/T++P2Jub
5XlAzEWrEv+9Re/xLUYNQflRrUubL4ShObUsgDqmQCXZM2bKtWyIUDTeILQfHtYWOsBGPr509QZE
tZ4z+fIBgMURNk3eFELtP7Zq+X9OD++ky/FdR9sOMVRGWKXDYh9Ze73tJlE9uUSJMVoc8lCoc9vv
dQ8u2I/t7cNGSNoLT2HKroq+KrjhQKdo9bnwj6lh9Fs2m7tiXYSKsCNVXBEpb8fmtdJ4Wrghc6eL
OoP8vA9g++GeZqNYDLtZDF67vb8QWnuQs8FPhcCPKN2I34zfZVV61siy5VkkPAtXv7uDZ1YxqbrW
54SkcGeC4kv4v0M8GKtI7q2A48nNfH54FF0AiJm6YQLDet+MSt18dDE4SS7+UrM9x/1BxZbGBtyp
pJ7RcewTvuolyhR5bqQdZqohZO29VrFZlG3Xnq41gNDESFu5XCbNywclLvqA5Y5EZFB+6YKiUynB
4FvGn6y2UL/W1kBzdM+8hmqvqveukFK4+qyg1b1g5vkz+X3zPfRpIoIkRtm0pGZz+hu/NNGtrsxs
t+5ZqAnl1nYtzp0hNWX/LFePjTp3n3Ft/uF6V+V0wK0vpiOFiDSwIfjZK3JastJSiaX6Gc+CcEru
isdOt+mrp94g6UFNs6eRo0TMRmQ033NPUFElzkc3f6zL1j2JoWF6tNgr+vAIMc9yo4oVlMRrSrQW
69xDz/eijRAk1QcSCq6FHmjp2kODetHTvDWIsLInOXeKdKVPVHUrHJhAczxH1AE9botz2iGNcPam
npJetD+YEVgNfqxbCKwgk6YMq2So3QmZp2cHkxYZ6kv5Xs0imUFrhtvbCEWwfPtrY1tS9GhVOEiu
rQsC02Lqeetg71V7YpE56Idanh6Mg4/u+qZW47uohs9U4UDKgu36YQjlC8QjsN6bFVpfmK18y6rZ
F0nmIL0N7UwbqFWXbVEq9grKnHGo58Mf2X4iO78Aa+MsSIihEckcB+AKNNgxB7Gfxqc0vkyOW1gl
jabyh3KOLE978PQKR9rkBm/LSK2hGhYfKPrssW5tXdODT1Cn0zUyFDbtJFt+encj9q35T6eLSoLA
OZJ4FcgvqNWOCW6lizkdqtiGoiN+cbdZ9Zqhmj7BcH+aRmmYOMVRdbAQ1pwmldXPCKac8lxK7wRq
SHXBDD6WG3SJGbDd0ubWsWJ1bfjjo7KOupmvcLkvbeFgqIIiwgLFqdZsMffLogSlbgtOQep48yHG
FQowBBxP78Owhkdl42PWG0WBAi1onLz2G7DwB835wy9/38/ekTj0FPHwMZ4mExD5YbBLJjO6FV3a
4wfCo0QNBbwBiGf5371GCPyuyFxMaz/GZB5kMw9tp6PesaPI5dXiVd4ftF2ZYPl4Z9Kl0yDvxLkw
rRubdT+JQFqt7DZPElvAyzpZsgUsHFsdp2T5JNOATcRy4lGeNZuLm/nOzJpwwLRhJgH/OYT9i1nk
igtZb7CsJ26pcFb2rpZtojfcEqDqilW8BpMHpLJbaovKDNKxUM4VVcWtm4BgE1tpLBfEXO9R/Qj4
7JEkhkOykOa3hXBqcfkArwnyIG9OXix3UcFfbhG4qLa1IOIxdcOEkO0JAawPYglTW59JhFJuEz5O
A62zfVoHU+pTRAee7/vwLV3yiEsOrtCq7muo1LYCkZtvchbp+E5MrX2yuKv9S8MYLkILU0P3qyZh
xTzfYgnecgbb4lu52v0heGKd8y9ctZFgROzGqxwl2rELOc85h1YWSTsNts1vHZ0O0w39uWve46jm
Q1CmGHt5uhVhP1b3T9Hhg+6nbhDGN3qZ4LpnrxYw6VQrB+U0ZB7O/E91ewD4bryd/TZNa2dqJRgQ
fiIked86jN5rrriN2LdlSwl4sIKNMBSr2feGsdm1LrTz4DV9/l2sW+pDobfkX2lCHvAwx7toCnCI
5BawUL5O9SyWDyMw0Qm93oNID3ENQA7zqWiStAGGvzAt0wq/wrA1a5kJUqSOEmJLKtO4Sq7ElX8s
lbJNHVUOsmNSGoYW/vxKu6ykrMtgvwnuugLEcQE2e5ozs155JW3LyE4Hpz8EKYkEFPgEisMMdNpl
/QE+T1nmel0oH6c5xMvi3XzdcA53fyjBfwXp/YJbhx0PfWLaUqkPbYORNNSjzE1eXnk/JlLiet0N
vfF+EpZhkZYp1RUATPMUVh13ZIqSnpf2j/evrSzU1bgaLrqjfhX3mkaVFMns7t9obl1OSowbWkjU
Q5sg1bPptN5HS6+qtAcIat2ai38QazuEl1pJ53wOlPvvCKweSlItQBFgAvL/KCXjFw+PjYwP4nnI
8A1A5jQIgttyOv/grZGPAwpghb+SvnVCXpA6D5Zjdpxd9cfvCsGlewslaNmbxYOsCUvCGaYQF3EA
C1Vs1puGd91/nWzJwL+JL36HpKOS3h2reOt9zac0iQ8JSUlxl81gJqImSm/Wtz/EWvJOqn4+gaf8
CVQvuPH01/UT1HcQW8UyZn2wT83gZHprR2aN4GJnP5VmT1YNeqN930dN/+sXv8XIgPgLt0H3HRX/
Z2HoeDPE7WYR0CJrkiW8bXPuVesltgsVfkjCNp1FTtAKHRspzCOxgauPQBCKl+GTGtEEMzlWw9fY
C5k3U76Xo+CC0sHTtp1VIF6cCY7wQ+VzhqmKl3y9W8Hm/L2lsBIz8cXBT7T5ftRAPMuzZq1F2VNo
ChBZh9NHghiuKCR6JDaO+FIYdcaZfzfYQj20OnQBVPVvlvbcXBIdA18QE5JjaH4wYyfOfiajfVou
4SNMt8q4t6Bdps0SmrIdHjHzuRR4WmB4tY4ZUJyUNviO+RnK708NhoxqBR77MHc1N2InM4dJ/2wG
LA0de8FhKXOQh7qpMu1sICti2HP9zQCDUMIEqBivmk44/aYTIwXs/hRQhFFtzMzXiPC+D4547/uQ
4eIrYe8XoKZpIjNuPMTOR2jJsVy4GhHvXiJl+yExavFq7MWzB881aP2DNEIUksgLSqUwZ4vKjKzl
SNkgZnSPGWAqVnPL4OEvXAzI+8gPSoJBKeuc0nRqkDRl+okMHO5i3Ze+mODtygMK+6MSSz4wIhT4
C+0IGPT6KBIyIU8/SRI6pDt94rJ1KNBY1Za0ppCLssAMk1PuQqEE+rahp0eXgrBXqXcO/D+wusd9
E4K+hO/yLhciQ+C6wDLkhsHfF859xJR0qYk214lT37Ph59HcdSyJIeDqHYJTQlsWc+lSTUB9+bYI
AIkkr5RHHgWVK/DScj2zBBz2YyRMsmjnS7VULEhWEVKDcB+RFoHmU3VTKzSeqy5YA5HIYpVPFig6
4WCIVSi+62mzFuxNBpboRLjMDaSdCoKIa7eEw6RqLC7UqM7/osUkoB4EL7jUMzkB+AuKq/KB1BTV
yTl2TOyW0cZ0UO0O3DdwKZd7wEncfHPi6gfPLL/lDi8wWEktQ4cvNwRQu+J/dUtiF7GCKdcevFKb
5nZk2OaqRsX+Uro1nC0xfQKAHERTwLHS58yHpVCg4tNixki/iUwEG9AVfzaT52EenJY2hzoI94hR
FXET2S32Qa+KS9rMAUA7fgJ2LChC5z1jsUByH0N9xjYeecjnbYf29dMgMCRIo8ApvSqzZuXJ8bD9
m58zRuXocRb00/fn0/vHnwhtYJajVv6UzmgwOErH8E2BfN+cGQH1J0mmaijlDgMrynt881ZDp7AV
6zkgF8kdpLJqUroofYNQ3FvDGrJ00xs4WxhZ5DxzmVHjUwhqHutFhFpFENNxzQm/jDKM3+DvzPii
cDbNHFHK8gRRBGNpf86M3oy0XrXku3QaiB/ds0GNmRwGbdkyimXLUVf8sdFM1OR0r531SSb0AenW
cj3oXpgrLagdMJomJ3xz27jKgq0eUnnlmjxxixWXq/PDxN39swnxs6m8oGUzKpXpBDc7e5id8B1s
7+tUh/rPf/DgMm+u/xNu1A/z7cM5lLaRj7++sJOSac1rzKCHcxGWFIO/CUw3gbvoWUhq9BzKuU0E
tELL3B9QBIKR6Jg8e+HZ+1eALuM5gHk0KDRqpj7ozG5l4sfOfLd0HMK64I4l7VzRWqwMbH7mq2vU
ouxTaw7U43L5DfqBBf7zpzqjpVsqQPYefH7Z90s1ANgdAFNMxKB0ag3RNJqREcmxDkIXVjWrD4q/
03feOxj1XsrlFe+AmVZhJGh/RTtf+Mv+jz/kp2r2llqQTEvxJvGCUYtXOGAKiBRHZk+1h0TbcAr3
JalQAf292kb/wFObw7xNgv/fnQ/xOrsRbzIc7AoNg/u0y+B+o+qtRLDETfmJM62wMqsyj3UaOQEZ
/L5GPypkKmgRwPyCr8cYSUqNAofa+tCn9yQ6oaA2QjRK79l753wRskY+cu0N1wSdKXLQRVvExish
hPuIRRDc8tDABFjNfamQy3QNzG8nLev19gQYYM55A9ag+Fd7ocbcQUVoIYLGYB1gljMaQGi4WjIF
bkzeIId7qh5QnRMVzKlrdVVc5XjreXaBQ46QRjQodr1Ea8K5lDxnIU8l9DaOZWWIeBJoGuLlKr+3
/cyx/tDmZ6pCvKAygJQA4C/gW2QOHF6EpwgWWAS/62BO7F33YF/w1fINSxZCuhqkVvQFh2TrBbN4
DPX4oDK4YzL5u9Zls0hoyCWw9eBGJUazmMZ+zZy4lVutxkHRtC7HoEW3xGm4uRmk0c47omgDHYV9
hduaFEVnF7DX6Q//yy3WaEgBeK325GLwDB/Vi3GEvk9exSuzSj7NSLZ5aRSg3pk8JI9MMy4IBjHr
gcO/Iuwu6tD1kvfyMlBEfj77SKxkxuwAZPd/Xx0ly5+p3YkS2pnniO4smGHlyAIHiZCY2l2jeRKp
yosXelrN9udbhe3ugLP4VAxW/F5Uva3hemEQ3aiCpk9XZaOxGbEU6BDIaP+wCAkhGYz5c+tqc2BC
OhRnAopNG+Yv1A2/al5WThk9AfjEiPvnlcEzZjvc5s1/Vn8qOc/WTm9cCD++zcOukB5n/E/yhU7O
sbGVsFHa//9kJ/GzgPsbqvK6EOGumAxG3+nFKLdhj7ykU07kpJz6pj8pS0NdK/rju1ttOFC6sVun
kEjrgo08LLjHUm9WpCUZPxr6lu5XXO8LbQvLbDBC2GPB7shrIjetIHdh8NQXo+RDLSBLDnsJazxI
7G8+uUL6c6OrPpPTlwCvPL8TxDyo+mMFl8QI45d0UgeAyrXU7f+qkBISdSZuiwsVoAf/NVxeGBSk
8mtqx21XzS+zBYIArHF1CjxY9i2w2knjSBBolOOk5e6SGq/aeP4C4rPLRxlCBLcE4tsb5OaX88M+
GJ7OAoDkn3vPCmokr6kV9BXN+TZ/GOzs3gI3dQKQG6ygNt38V2PNH2OAovrZ0ylLzcIfn8emITwR
xuNC0ejcXnydyS8105F89ySOg8O7xOf70sfQxbpUZj57S6M3JL9YadHgFAMGYySjbVZrg49Ri4CL
frv4+fGZDtHvkRfvsaJCG8wIMgLH48trh2kiyYdJ2X24V8IzRQSabpIvIt3w3ZLZlf7uIWELHgzO
6XwV0u/5BxQZUCHYgZeUmRpfS1MLxPsgOUEE4mRAbCAnW1G/kNdnFwdGco6CTonMlQfI/JeOcZsv
oRgmeKIyFQTqZTsSU9x4GFnId7pkN0te5zgL0+LLcvKrv+8JkNr/VSEf5gM5EMxBvEs6jGD1lsYv
0BDtYwC+Ncq4LmO8VYhSRDwvgP7ENC3Q/Qr7v0pqfkYnsUvI+gLeJ/k3oG1a+sUcrvZihtriEFPH
fJqnmMo2zUZfiCUnXSjA7ypuRFXg3L1f5pUy7di98wgQ/Psej/2xBi+QnGWRH1st+DuHWhqKMTOA
5YJYTA9e1Bqd1NTIqsZ/B+45BHHKMWtPEdC97yMkcjI4MV6+Dk8uBdQp8l2oYQD3utiQ8jG20qgi
hQpsqWM/JHSObCfvlyGZZ4xHX8L3pRzM4lGZASz1dVBhgpUeBi/EB/QuEhkkYEbpd4O58BJ1ZMc0
iGUQpeNVyw8ZTZ+Mnry2Co1cr+kmLKc5riAY6u4dqkVXM1b7ogbgi9IckN5X3kM0nxUcvwWfle+s
zOGq7NOVCGY/OB8GfkBrGAWKsXhXBamBWTegmopLPhxqCAsqudkLAf0VlOLa0x6AVMtnMBbSKvXz
9emn+mdRMicu8vHAzaSeHM+MpIppXwYhguSnEd1PmCBaAW9DppGXfqP7mWM/YVGxt8ZEQOc6OxrX
VDRZF1/fwsVCYzOjNhs1b5lrfuDkEc9wcSJDGNMkKa2YdfCHYcQ1oft6bpYvPIETww1UKmQFryG+
RZOmdS7Y1NZVUlmrAnRHbODsR6afJ8ZizR0q3gT4HidaIGP9aJsFg6ucc7o4um7SEbYZqxwQ40jZ
SrzRbl+Y4La0gChJyMlygLW0Yu2AQ2ljFjX1pISD96gVUGBmhASOcRGSZ7p/VLWttJgD6h/pfR9+
FrN+0f08faazmGrXlCjjspFFGojBImFofd2j+bV5PgE0hexZhpysqpSCBtp+Yp4jQWvouAMAxEiW
xPgv3OJ/RAH0EvTF989XlGdpEhBlUqIR2zTzOQjqlZtU48HWSXP52cbGIjXWdCkbkzfuDhMjf530
U9PK+HmDszKXb+rFGPs4ttuA1xLZ6TkGGWROqrcjFbDM27w4+fySiRWF5kO5aZycjdIeaUu8BdBM
peZShvdHpCjPZEHtYOmhbviaVKRwnAWnlD52Zbi4wH0nQyuYEofeZ9NMZOdn+Rf8QT++TLmj3nU0
mFwuwEwrjJ3gybY8bSGD+Wl3NUd8vNBfUwBQeY7gKX66Yjcy7awgfNBDkfiQjJbe6+rgfoflTj6v
mvcx/e2ET1a6iOZv01ZHjSQ0niwr9KUlpLwhpdeYIlg25/pNc0g86Z/acJofZh2mIYtxh1+/QR+s
0RZNHw4s3eM2ACO2rYHAypLn/6zIbPEvUP90tklg6vabZUsIir8niP4vHzWTILDMGGQ6JpE0UInG
BsDaXQyHrXVp7975Egto718ELLtgRBEPNnlV1/h8pj3MS4LSLfYlmCK/mPtdIJ7XGimivJseapRN
4TyWGKt+n55SBOGod6QJCHZCZRDh1gpaZj1W72NB15oDeDsIUVdbzZbZD3ZDvPtxF2eCrbWiF3XD
MrQNCdw8ANDUE9cPId6F68k46qTOXrcfcIF64icS64K5YEqpLY+asKQh+3VlXCXzvKH8R7OrjcZn
RBBVnzAhtN8SzugfADkjEzjNocW28/N5Eqndz0zRbT1TOK5L/P4Pqoum5vMkU8oLLaots5AdG2O3
sXcu260uI7NVY10h6IA5yICs7GQXOUrmPHY5drARPge3BBjnLd8oexIkuSy2uNazpwoHkoOXXhxn
+IxRfNpXSfqhmtMpOcwmpJ0ZEiAi16dmsYsOLnc/IRdJX34++5oWgNrVbY+OMJWi3lWjBEQqARDl
l6oqV8cfgyijzSHYhmxLPbzhtKAnxCCenMIIVyNiKEAOyVELKJJ+CS4IexJznU2jO36EIvrHhji3
X4UJpMPmxQnA7ByaO4ACUxhM6rhtcN3JKqyqOGMwmeAxeDAB5Ka8nK0jBScFwkTpQPlhdZNieeti
v/i6o3swWcB60JC+aC/BNPY3uuXlACIi6lHOSfbYRwTxbzGPKpqgB7ClBw1kciX6PjCIzvPjWZ1B
rGMMV/LYHgxt6KNRGaLokQkJ44MdrlFTo4rZouI8IKPeT2gAPdAYKdpKglHK1g2f5cxY9c4Nz1hr
7JV1hmSCZrJJhVuVENwTbNA/2pdaj30NWtvY01TuvwTeK7xJj0gz9kv7oBYKbMNkHjFK3S6dSHx5
VbJVZr//ZYd2VtTleIagleQWGtF0e406A2f5IDbsR0U2wiunIzerr/XkfKewlWW7lukszfTCtGxq
/5reHrI5dp2YHlDyTl6Z51tm2CPuQOEh3L0VCQEAuzzK2/KerHjj9nopQIcJVCwybBDSGlfdQaPp
PJ830/Kw/NMG5S3G/acnMlSXGwMm8RQYrjNryg1UfRTZkSTRiu1WF7KKnFaHdxc8O70NfH+ZDNXh
Z3fGtC35ZU5sPYQlpdr5uP4V3clKVVHTOWc0/3TVh8Pk0N+hHHfBPYzxIJCDQCeKuCqs5ZQrK4+4
Ww8wxsQ87MergqrlGv/B08OQfFaz3ZkP/iA2iPzZLqIdmuLwK8vxwPtqjHXdBtiSSJfLtBOcq89a
r+jdOJVtZFp/Vj70Eb0Dhz/1l1pbMkGyPZjHKQPSepmCqmcGWLBtPLknM6AdyQqReDhC4QXE0lDu
85pz7mHuWLkjVBA65nVsG7Rw+6tOoONvoSaSA8v8gec5cX1dPRYnaVlwjCJGe+h83hqnuetDZKfn
A+9qf/6n/FU0zlPN0gwM90As76IE+cTO3mbyxoFFwSmYaLqpwIvjLREQkglvAQM8cKNu82lunOEb
/85evbaqdp6m2J1D85CWgP3sODggQjNIephsLFTued01g5aJmRoU71ICBCVOVhf7DZEqhoZ+Y+/i
+OES9kqZundlizI4EK5neB1PIhn4kF7W3GQ75cOozLqECrGfWe6r1xyz4d4cDqZlm/e+31xq0lEp
UaSvvhqz36i7+y+mjGvazRjPRBfyv1r53Y3fCwLfY+46h+UNaA0Ne5vgfvNCDrPP3OoLdXEhdNq5
CvtJprNDxYLufYgzG6wZlhw0w7gnu6w9s6BTHlc31OdS0tf+TDKSd48xaa+QnSPwSGBVNlnLjQUQ
T88CLFv33YUlYr6WG0VTUOi2e5pIAWEHX0deRjibHxX+b9PCgMo8QtZ6GXuExJq4f25R8GOwHmMV
zeEjQ/B1swfJVXrhsDAc3c1/5I0fHPqql5VDuArIutWxZ1zp/XDL9NeZ3dzaG4VVKKoFg6UTj0ob
pd2+t6x6CI9ESp5CljST1OjVcosNBsjnGy11Zmyymy0ODb7Y2IlH49rm1CJ6ER2Z16XL+W2n8Lul
3r20zvyAUuy+r/zldHrbLTG+SfcTnLyH6UO+rZHU5GvynvEMWJZ5wzxa3lvL0G4K+xJ1B5HQ3MrL
Nmf5Hhog8eBbcZTByyJBKPQagvvUX24+LHO7bZKi+Jk5NSqDZL/gtY9stiLBdsN3dPlvQptBvvcq
qdV/huIpl0uoQkekweyFJ03TzrNHHyNG8MkB6WJ7UuKKJK2aZALDCIzuOWkJgvW3vdKPnoO165D/
9x9K8IHq6sKN+0zC5H2h2NqOIUkXX+2HTpvQAHsU8mqh66mP/FLXpcIj/vwCLK4VX8vPqGTz5xWI
K54Y3tEjdAW/m07/sUrmZ+zVvw1n0WY+PmDK6XIqxILIAQCAdYt8QDDy6mRr+7BRe382J/57BeFt
g2KGdraKKe623lZuJWyHP5OU6h7tYK9sO++LW0588psz/UBiMjj5Wp0bPuAqqs9IoKjqmxBXCXZp
pMwKTlbVjUDNrLjKr5TvhyxUXaqqtYN62ifpk+CoF5tKeWAXZ8NN+zcpdpbNWtDNbMPmg1Qhbhc6
Ov9HnNIGMPwr8wV0dbwVu3wFpYgGSHTrNTVeWexSD/AssZUf1zBEnv74yozRXbopoVXuWnuhgSMa
TNHg6u6poIOlJOlfHE0ZM/X5pYIEcoqmy6sZcKl7f5btF8DB7VU8NaP3sP4JdcGCRv4FDUm1Ik4l
WoQYYmxIIL02UDvDYldcu7UUjVgdfa8PNj2CqE58hdmKnqJ+D61ghmjOvPlXxHnpdhIu5PM6Zw7q
68qYtZdDLSLGxea+Gs3v57V+iFOunbrwPlVzTKnzD0zL42zgR26tiZGIIHADwsgwR0LLKnrzH3G1
7ZZCKWdp9VjAvQZsj30Ykf/wT6ZeAUCHorJ6iYtmOnsjvvXnjZ0qtckYOqWJp8xSuNeHkOIG3VN0
fVrIIV/yEsy9WNy3bIZ/on8EwDW0g2bu/zHRkNMYNehTbY1KGq02KbVSKH7Uy+aO8rIicaVSSje/
nR4kD3Dlol16O3z+K/ZdQIOeZ4Z65NxLtiK23DuD29FeYDDD8yYIsLYt7N47pcWXRi08tGpVlQCt
SUXcT2K6vaB9UWqHll6gJYOQhrOOhaElpBXGDmYdgFlUg+mPmAzkTwcI9nLkbP8OJU2YKdSnA3xF
uLy2vBe+GrFf7/32gKCWQs9kMlaJEDlUjCH496MvP/u5VErU0SR4YEX0ZZ6GT1JQDRqrYNR/y2An
6PsumT8G3cQw8cz4aZVraemomvDkURMSU7CEsn81GaAkdjezRSKWU3hmbZATXSmEW09bLvKhYboA
/KdLE913iIlr6TBMsuq7ziDaS1gkBnn77vtWHYIm61cho3wPHYX38pNwyxhl3zaBtxmYtKCmz+Em
Npdlc8WdqILHoTIfCjhep4TFKE3lulul/xM/8pw9L1RGeRk6LEdnByDq/Cbht+MhaHWDqW3mKCpR
hNwnjvPsqj1hbGw7nX5hiQnENBQ05kAYszflTLLHrGWNzWRRmeRXaccHZn1ZJKx4aUPhB9+6kdIK
yBc7jzOO7ejxlk/VklFLx47xAZ7TdmdPtHmSx5Wglw4NDw/FSwmuiW6UWGnHztXCT1Kx8PRXb4bV
pRszO6xGIYaMLIY2bewIE4hmpeaXhZBQq0eYRzKfS2sJXPUbt9+PkaRe+ZmZhqSCnd2RbimZQI37
zOalNz2Q4y5ozWnEKge5lOgtfC1K/sFKXvgsaKMOfgx6mfabm2+fct93RJbxQcSpqWFHxu81Zjeg
EpVmuXXx8f0ZCgWh7tkk6AuyKM1eil/9B3BJcjAjJYxa4oxMbNayp/t/0vOijdFRcgQANHTN7pZI
xI89EZmica7z8UPb5i+tFBSv6p2ZkUY6aM0zt7n+GFKiU0LyQUeBzRN7uV2FfQJh9Ng1MGAays+8
h80xA3nHCeJvMUcXcLxlQ4nYzFJTJZf0lqxwnSa2IFc0Si16iyw2lpxcMaDNYIobwWkery0PnfVl
e10hWZTKy7RVCITRcRnyc5f5d/0qVAgWccu2fibNu5UXmM53rgriUStwmxS6eRWIHPgAlGcdGL5Q
vHI5v0mbnio4LbHiS4NspCS8EA0ifBU4PPXI/eOLs6345+7XGu/anAS+Ow17qB6uImhRMfGXtUdN
ZWC5lahSNaObYO1mkMbW8SSw7Kx3fbvB/jl5W1vSmTA11JWk9oBtHx3V3kCQTtyhtlqGCm3W9ACk
S24ND0CCT/UkZuaDuppBviS0HN9xhnkK2eltRkmR5Fo6nEk2dvWH/fKJrcZVNj4sVHlTRpyY5IG2
4ejnpA5CgWUm543xKoY5JAw7aBC5mPDskDkCXENHkpMG962BLSYi6qQ8HhshM8TfXBbUBZqZgAR1
bfMln2Ilhh4WJ89EoDCsRcQaLJ5NR1JedLtNwZfZg7IMhVEH2AKFE9Tux5qpWDZEV6n+PJcbEVOY
ZKwKELD+FA5LOCjzX7iSGn9PvnoNFhiw5Ss4WbliK9Q+0DztfxXL2zWW7JD6cNAo8XgkwW11wfO2
uKQbipWVkwC9z053JgLk88st5yz7EvSGI6ACaHgsT0f9dqMRMgzqYNxqDFK7c8EHH7a34cLXJC6S
xfr+erdJWt6gnL51iwYEiCct0pTgZs1aidduWtmGQHrLiGRlaA57bZIz9YjVuwDEUdIFuMq4yPEg
3csl2p3Chw9aAE6iIgOl+KyV86yeJX78GLp0fKSzXy/StZZ0f8z/cEfw2Ox8u4Qu+WoNeezL3Qdm
iJU8ge4n5zxtqZ/nbGph7tSUlDGoQf4Jr4oa0tTzt4pyUIaDmrJD5uYtY0Dtqbnxd2gylhr4pB1R
shwpwKVN4sGAaWM96EYYaQKKd2gYGFSQ0vZBOk9Pp5ntseZlxThuzyjEzUbDsgymZZ5UXmPu/kVc
FJEUAJMADGdSoTVTyHrNxL+/NYhV9Fr1CG+yaW++uw04OzEYxGJT6jWdj+2YH6T1NmngYc51P3O4
IjhbRDN4hwIpLqSedzEMvQk3o1ej3bOUCjpKROpIBNJHlZtHp281fXnHop6hnDNFrNxiK8K8CYoz
o9vQpmYk6ogbJOQyQYS2Bute3itH5PdEoedZdGs/fKzsygvkWeAQzXd2pVBcHTlZ+bHf/dGDr8JT
7shmdYcMmN+7TEKjYzkoj/2k8cj4Id0Vn3IuWIJKVMejcXi7NW95pVBw3HAw1nigV7cCSoMvqBV9
NpoQdSHY9djxf/+3ZtoiKCah6Imrj3Ut2KPXBLyv+N7sQpZ9x/8e8GFTPW6TXXAjvgCDEbwm31ES
NAGAikKnLwt2RI6I0r2unouPPs+U0CRrgrBQVnYNaMkNJr9yRqHjRglHlREsd6jfR0z/I6ynOrjr
oAK4w3q5kkM8Ge+FlZAmflnnfFpAnGy9IL4USl75HxJasahIsBFYqRoHoPFgjXh1fGcUF/sZMxLq
o6tvLvS7WeGT0Z1WW7+bGKje3HCgpkgMEL21eCwPgx34vbImcRvGM3DGlFdImQ/Qne2CIIWfhasS
Q+dsJypI2dKV0kdxjmY0X8KVrqLzrX10qoBU1DSdLTTHvgXCR9ljaNuLIS9UskB0/s6+fDfvTPDN
DOSR3Dygaos8C4VWHLeXA0RROmoVlRA/tAJV3JXR7/uW8oT3+qw6lISJSPEJcumpEqSTSxofJtrf
IRvB1s5UvWB+DLLauTUmLTvVwWtCpA2nXNs3t1HE1tP7Wrt2U8t+H0yLQgvwg15KKB+z8VJ6lsW9
zAHAIDeQ1ZSDziCVX7fUgIJqGdXY329MN5t9n4P+Me//CEFHZzbzA57Jxe3bIYUlusqBTkzQgSE0
ixvCp9ANt8anBbFE4c/0ijql3mqjXSlOTmSmNBTWLKXAbSTn8iKrYML30qeOgcP4l/pPNUcLfX11
k89QYtOTlLCIHs7iI+DHJl/Fr9Cp/t/L9Ra2chaMviLItjkvAgGwv1rpdLTi00ffrpSzbeLMJOph
wa/A2oSTT7JXXbuN5gUs1NWPh3QALWMAF52pQLmv+xl5jTGwz05waOeBEIDq6083QOCIGamiIjXr
F6IoFS00gcqWpj4X9R4o1BFhBr5weXtVindsyp4u3FZFNLkmvjV9qie+U/70DbdbrpCeKxPsSBrP
uzt6RLALI2HJZ/ocHq3/b1uZprsTt6xrqYt2JJqCT+k1b0HjPyc5V0H0kVK6jwTsPFWhRNYhHE0J
nleSb5pvM9lRYVyE9kWHEDryopI8C4LXuwg1b8seqrnHtFOqlPvJ3RYDs6Ak05ZdPnESKQsZs9/y
2DTXBhS7AP03Q+nXT00OpWRpB3frvpvxse4jVSAI6DupZxIIhGgs5rtDVykmQPhFrBTmt2fbWI0c
mnZEkcCqEdmvp6r6svWe5KgcYOl5CcTBKsVVtDHi8mWAE1BKTWGPihyVBjHf6MBIEMWWW0vALKlp
8zL4k/fp2GgfYaU+3xw4mx5mQigYg0+5Q7dSBfIceLii0+UMEWCoO63MbcdUV+2iOyPhFAWHbB4Q
1XZUgM+HBy2gxYwwrD0Kf2En+Fj17+i8/JkOn4/cJG3TZYKq6OlK2C2+CFmsEJDdYfN81n7uMHcu
rklnAQ4HmUKfYksfz8po9IRkUHbO83/qzUn69nATmYkzoiZM5TYrD64/KyZmalyufRgdWBmLFqz7
G+M7WPljeQPf0b3QMhJgaEGP87EsEFq373kWWeNEsWL1twyJDkPQLn9IAf77W44zI/wanB2aupXt
q1XwrDOL4Moh3jZk2Wilmq+lCaH56rhIMUuhBQ3K0nFSGnD0KVi0UQ8HEanMJx2xn/pPADaAzICa
wB6QKkw+HdP3E2l3Pa3q9Y5O6uDnBwJ4eWqCXYCLIvhT2tZewD4uMnyh41Zgx1cemdRpecxEhhNf
bE9uLGtHAzSr/zQm5rSW8vThVBCjhEE1tpvjNsW083gjcB87+Mxq17pyt6sE9rEyq3H+m+saxaiq
zSOcUBWAklx8ib6FFrd+f2CEJz/Zh6sT3bDpzuC+y8Lu12V8Eg6TdCWTEtkXNw2qV99C3lGF6pMZ
8awo5uqv0E2JIGq5rmsO+bSzbh0ZD9bNg73D8PQ9eoQ3JgcZkZ0cOHoI0INnBlpcr0hsk/LTJ2ci
N4IPk5g97EVcz3/9M11EYk9bDagNzdUCfZqdpuquR4+6XzW8BtsffMGqdb93TLTjSakncgATVu6v
yaDc8DDSojGb+4T9jefABq7R5BG7IvelgnXeDm8BnHVqFnLco1WUWc+Qa9hd1Lme1oGckHgbkgov
H3s+vuSvt7D7eren/v3h/ThTWG6obxy7QrpH5EYHayeoe63CeGwPhGMBc6Join5J8xkGP5Pq9LUz
VMiUIzFtw5WhbCKnYPdVFPNPfMQStv8A1zxrE8mBHibnnEIz6AXTI+9Oao7lz/vzrcuZYorsDz1n
XRK49L98GLCp8ZKaqaX0IWAOyGQcUg0oFzGuQeA8bLcSGdFKZZ2VxmPTnGI1Vd2Ex9Gp4danzv7Z
NJ8dMjzNuKEepMmtPy9CmeWbINBmOEvmErBbPBpACZA1YAPQxgm4EJTMRZp44eo7IUDLt4jr9wI8
PXWB4k7osP/i//bM4OcokPF9BQ3VKD+nAEdlNpwXo68LFrb8MPv5h9eKq0otrgfHYtk8AlGlLznC
v2Jq3cs5mGkRAp2MI1HFOHGoCQYsZWurTQZ0/qUWw898GvnQ+xx18oiB2a/zC1kouVixYuoCo/6u
ER0+F0/41oa4Ir3HRg0prLrS/bkwxEncBYIUSRnfnvO4167wGUTNWFqj48bJqPG22NDhs+88SQve
BmdRBN5JJgblR2FJm2xiyc6yxOVDgnAAfBSrVGpMslx0aXFeua3e6o1gFhSnfB2EsSuwrqFaok8g
4TaEUH8/nCqQXaL/kQkp86dS3M/wldLunGGyziOExp0h4c2YKruOAXpKO6KpiEU0LgBJzM4/fwZt
OaZlgBmIjlW7RChgReCjlekTy5kneudGMfUao/uHuFQWwFD9aAWdGBqJb+PiwNp9u4jbabFSu7+R
hgZjI8341Ymx4mVooWB6xRDKQIIQ5/Yq8A6UXzg9ZZmLnHa7eLV48kNVqYo92c8/8ZeaHkXn4WhW
fctC5ckgZfcMG1jYiJbxX8Zeb23m97p1bc4J1EB6QZoX9TeKn9eNJDp2bHCxZONZXONl5DKPOYHb
/QCHgaaDfT9i3vqngqUjp4yUF8weutaJkN76E62V9Rf8nGKSn2J0Nb3bzQ2e2wvob0h/NdtEl42t
Qt757dNnUBHizLTSo+tzx7ErOiLJL6qNP8euq02CB5iIBe8wAYYWhkiP5mWjRI3hjNks3S+AnHh4
8D5xh/2aarvt929KSqe8FEk0p0K4BqjBzCfM4TZ1rmXAUoLExI3fauZlaMVBLaTE0Kb7opGLwIf8
66nVii1egeVdngQmJIEoxKGh5jYYOfNLqZmrUwESd+W0hfSs6ZzyYu28ox91PB7E7951G3UnGZsv
Xj5EGyYqc//4GcN2T9wiOzknIu8WlCJSSr2AJHAydegJuanAy7D259csZv3x8xRIxutd7a3jWT9F
BYVtuUiARg3DI2JdBRLEOACcYK0bbqHjNPSty20LzxeI8nHUYB5QegFRT329a179bebJgYDu+Gvn
oJV5aNu67G1Km+yGvoBVUOUfieni34eHqgDqMYKSTDfhRPerlAhN7ml8TRPgpZ/PUd0IPjyo1NiC
1wGsY3+qYrwNCK/D7Y6mLiZ4OtXCy7E9ZTQI0NVoBSnzejvwwt5HMOCejtBAyjY9vW6v163Rz8CT
xWRv3A+szVpujYtOVNSLEKafHxySbO9Bmw5/I00x2f5plqT3yVv8g4Sgzy3Hu/qU/8uOSKYAYTCl
ZeIHQiGRcDEzzVsYxjQosPoKClEPBFZ02hvUNGnQ+wAH+8LCt7NS2bMJVY6nKYt49nkZ5LRZL48D
ZdSOwNEXUCBNgbQCLdK2AjErGAHTiEqvzC+IUr0Cg7/YAhWSTVotCFc547RemjP/XqMjX8sTQzmz
QNeT/3wFFbxkd9S+c54Rrv3xHYBPzFUCq4VhqR37K7qhf7Xwx219bMSBeRaArZ3ofUEpCk262FJn
8QmX5sHs8zErLEdIOlwT9RKR0IdCrFkmy7Qkv1fubiiPkgpNhOMHqcfivxGbC9n6uQCdNkHuiKTB
rpGGEKWRhlwStj+njey3U3e9lCJIn1GPNsrpTqlGN60niTH/c4FB9XeGm9PPjS2ZoFL9pW/PUv2+
Anm1sb30ujpBCNfz9YvheEnDJL3/g2aXRYUmoUsjFFvmbbYAsSkor/DH8p/ZxoxKVyFRds+iSJai
AiaaeZTwWFPleRt2RWiITtNIjEF4Opxa5l9bsGH1jx7p3R1PUz3HxemXrjDTafaVTDsL3wzzS7+8
PpIm3o9jbiCB0vrIAffgy+TJGgBNCDQhRwnVOtzVei0iBqsOwelzeT1bd0rRTmQRLT2W2S7MjojA
X8uAlhcnSXPxAVywYpAg02O/23UX9wVoNocoBSZZUCtSm/2Qti7VdEI0SnEf9t8vE4prBe0AqPtg
OjWBb7rFFM9aSS+noFHEj0ZF+1mm6S0M2zjxGlC5ysijNffZmUJpb6CVdiruEFBf9+LX1h2YyzgU
h6w/ncbPgpMDqDRMkYGDmInpe93Ch2lsbFQeZlw2on2s/gnxfCW9hkO0dfmGaEcDn7paDJPIO1i6
4lce6+E78r/Ai1CdXJofVUrPWQmQ7qMSCOVdPrE4cEGoI/dlRykWsxBj/ipPWYUX2U5oWZjcC9+/
CLMSnWUPx6pPWtnm2adWM257VTLV3/Xveod7f9kW1Vvu7cFCqr2i62GJ17jQKB+UTEYxJTVtrH16
LGwSrXafjE/Zpk4jf3PXNdpQ5YsAwLf9dUh3rMTkXMWmNH9RYkF0+nRIz7mrqbuzEQPmlkbRAI+k
YWK2IVUUTUx/MH5+zR5oiRaCCee7y0Hb3o5FVC2Nlneh/jKiISnfEwSiy74zTXsEthzht/zISnCG
dSfPdxKErmDAO24zUhcMy1UQuVj1+O6lbCgo4g9kqsl6TCf/cUCU3HY5EKGGjnrFJ9pvTBVpVoZP
l0rE7Dyytk4nCZ1PBpGQl61WbkuLkvu7vCdG2rmSH+wtVSG2LxKucfmCVMeizlLvkRgaC8T0ec2T
q+ZILsPLCR3k+XxzMzpLIMQHHbLGWWT19A/WBLzHICTrRiqNb6aEn06zk4nlGMEjD+ZeSVZpyUQR
m35SjmdDj32W3UJTSOHwZ9SEQI4DhBAzbfl9S2B8YTmAztVDDsbWwBL+z/nKLpG0ItEE9epKIPZ+
1mYzzpRD8caXrZ6LQF2+hElM7OLCnJayVqhuDWUyV9dqwS6bq3mgXh2popMtvYp5xzUgiNc13hjT
3r2IaTRQ4ekL5dorq2P6Bzj99CTBBhTat6XaaAvK09gBd4xbu41NzNA8xPMKKTSTsp6AoFCvrzFJ
3XUdZHkDurxA9kaeirI97Fr13KdPyrmZNFrzaFmk82pbV8T0QJa1eT0/H9kJPhNpkUbxQJHgFAk3
2tLAYLr8Hl1KBDuIm/vDzWNnWqqNr54QtTH/o+Nv1yTWe34Vt6lh0bMHaXOqDj0xzaE6Z3dJRRHO
jLkxtBXFUhuRIx69mvWVumgmYZhPha6vlsZJx/zshBri4V3pE+PCAoy1NLJs19wlZYmwG9g2Zq+E
s/MiPqAMj/D5J5aoVWjfaQDtc/UEf5P6bShiKR89jctgUAnnqiN9DzzlJ0fXUuAbFqamGkbhvDMA
y38yxbXDlWYi3Tzuz5rvNZrJchx3jWlZtghPR9RlNpKTTvMCzKsiDGF8Co/xROkcl6MyUBXX+23L
7kNn7XxyZZYnzDV3lpgdJhnXJ6884RtmhN611VA8r5t0fKPF49z+naA+TW+PrS+cOvW9CpcE5ytD
9KyphVg+Vd9GKvsdsKWO6EIJEHRCcoXYNh0eGdi55QB4K4YKyvWilhCjNqRqWH/6JTcy3/S6T4CL
ZduxNqY9xUg9Sdti00/v2vOLUjpymeN6uuwr3u28Qxa6NmGYqxMbi7uMoULotDXPQ2FcbYaSvLn+
CayxqN3EyXApIPSZBHsVHIPqRLKqy+L41TGY70uQRCX9vN3mQVVFgJgliOevCQPx/wyd3kCnu0zo
Xt1RikWF0eLPIlqjmBblvXXKWa9EdQxCN/A0kZrZJF8FKysHIMrzvbPsTdvW5nmfzaLQyQhLB8GU
T5ItA+EPAIIFk5//jU5oWir2Zi8cGsMN0RWQ9Yq/wQvfzNVDBN4k5W4nYxRjP5AAoLg7/ReIqVjn
QhJJ+FDW3xtnr2oOh+jUeJlpKTzLinnE4ggHzk6q3n6Y3ILzC9UUF6cpQYtCsRKs8H2jPw1T9muE
E89xzOmhGIrwRTcUbRj3pKfi/GugJwSnuKDy5IuKP3fn3meoAcHJCSbvJlMHujJfEssQREZKCGvr
Fp2O5rYTDkypy3NkZtsBZl66qrZZ8WWjn7y7wZG4wSAfJW4zxmBhlhRQ9Wpw23E7jtQc8OlD1rih
mKJZoxGv0qB1CkAfQYEZ4GF3HApwMgVfQFUfgv35ORiRV7QJKN6g0SZqDMF8dbZHEBbDoe6uOX6d
wftG/OiEfS/WBPDXaH8w/AsnYoevbECLuGJ3xXzO2qyKfV0+ITBs56XI8rAG8E0QB3oeqGu948J/
m2QjgvPjvktCb4ov/GaPHSn0mAVKU1AO3FTn06aVXb2egktmTMXoAK/FIaYv0N1MzXglHeBzC3UM
k5FM8DNI4cUO5cn2R6mMdLLOPjOFt8vBBxAjaC4jg3wdz+GIFZ+2TP9+Vsajbw5MgQQQQ7ZDhCOX
/8cUI4/d87nJB6qqw3XYafSJjeOwqzBDAFsSZqcs/9w0THK7H1+A8wTfRR/CtUk8p/vy7NrLuiif
MWk0cq6Pt5ram9o4L0A9NW0xEGNtqfCanVx+FUz0dj6tfeoQbsABEp055/8nQctoDO9kJQCxnoBM
hF90H/E5TuBhXmbJ61YTaHpjS0KqXiMQR7ZVm0D+8NJ/jAhaGRaGEyY8hVZ0L+YM8xtKOr8UnEVU
CyivPd/lHcI9CepHiObvXFfKtgoa8PEqEAjiC0q9Qiour8ockCjeTS+ddZBGn4TO6lFMt2n60V2g
le7wi+7hwGcRoTHympfqPDiyBDy52gdPxijGCpUTQX5xBd/B92Mm2HDJDmFtk1Ea2GqOBwhxFkTd
4i0GPaJ74p9+fgd44ek+Ga2joTVjN3JevI/ybx8DtBio8eCJLBdUcqWigyZigJWZIj4FnLQCwKVi
4uM17JfsFEtmv7afYSICqCxcA65nqwzHT+H/fDb7qV6INbC6gdCTvmNBLQnW0iM9pv3ha2vabkTt
CugJc4/c5pRoqlPu77Mq3wc3CFIi5p/eMMDDaeRdgu1OWBinNOP4tM69f/AZ6MZ5YnKfTpfpM4PT
7yeCRsqK2hyLCxBfhVrq82wPvjDLUSdQyays6ZND/M1vbXyC5ZtoFPY9TYj3ebgMBz48thOIKP+7
W2wQR32wtV8UoNYzZjKT2/GhXDyeMPR2qU3hLvrKYApoZA+MdNeFSljhXBMSUwOwx5Sv9x5L8TZ/
neppKgeRkYQq/xiMTuhl+SFWlMwEdEhkbPhc1lb9FYltB9Fw7y9rePiTKVNfbdfrLq/kCJgOrFv/
RXMKlTpSWduNwgFbaKm30rBT3QDGbjyuN+wOq7+7jvP++c0bz7525WeAapmPrSwWB9iqyaRjHE2v
Be4KLaVCsKjqXx45TatL7XffXOLZLnuRSf6lMvRQ70RO6se4MCf0l4rcSnC0Ptr4PonNVeZTu0EP
1ORtLVwiVHjbSCx1RJ1ZGik9TVh4Jpd+zfxK84L+3zwDGmZr3Kr55Kw0b8hMj4vdfRILoZWoSbFh
hkgwd7Jp9HVupSJgCGjTD1Mecsljs0zJvX1PG3P+YGNGxsihy+FbMjM8aW0evJI0qbsxEsyx8X40
ReIoObxRQYXbc7c+/Jkth2r7BhBHZ6tSCDJN8tFj49wIpBOosGUQrxFURiAxhJSe+HcmijmcuJ2y
E/5U3zewro1pvBHAhFRae5BaUvyETXSKTYm+jsiaYJjpzj1N7WV1ev6n3JO0UbIRJ5+X+oYR+Kou
nLjGrWEVvX7vyY9HvHb+L/xmgiebNNJWoaZnl6Aj9Ksb9su329MiALPZ0Rq+1sLQBlhzsxpuSfQQ
H89ZjvTxQHz9/uZ78PLCE1c4TRqisHaRd3PHBZ+nbSWyvKuMDEvGggoSUGNTgB2CMe6smZAZSLnt
cHe04q43F8cz+6K7lR1g99U0igMAUSRe2cHkpeDe5LXlEMuxvUbGGPE5YqSCqYvSftC3wXtCh/r2
1/+HHiIOmgoN4Dr95pm7ZwpJXOTb2gwjOu0BFrCv1yG3zs/6/Yf8xXC3nG6pDdIIblxQi0OnUXqp
czFKciwqo4CB2+nmpbQX5ZSKm9Nuq5esF2inSpy7xs677Y5/zykgri1ZV8bMIcxenXkt3Q0WBWLF
JMJjY2smHs/M66LX4ktJWJji93edSvt/lZ5/xutvK1MfQc/3OqNoJ9+iXu89RPyJ765x6MuN5lB7
sfAPMGGsWVpBnwg6RL87VURJLdtsZWbFH2Xvgtxb3Lu4JyZtNoCDnCkNxtuCc8hWbJoLDPltZl6L
1KHJEy5MYT1pbFDInug5XYFkN3NKIOPaWcNq+0ZZaLTSYgalCnxMQy8KqYOzyEaW4kVXuVUFmopS
A1527StBG9BEI4MN33rW9W/jtG3aOQdtRIxA3WOPWsbvJP5r26YaTiMqvg83eslFoch5ovZaAiV/
ekvh0cGNZWv/hBJetqxazx2YiTxgWFix4MaHZxP2xskCeiY0LsU9o38t/2vjCUDiPROkdnXoT7v9
eiAH7YBJg0ai2Z9cTZMFu2xpPX2kBOsAf5ujCtczi3Aq/kWg2WwoumgpbCe2pP9vWbQpBOYormJu
SK6O0O9Ep7iuSIXlxnUdjJwyhixE0feXLjEcYyF8TBA58fPeomjXp7bSEnlA12FvGbv8la/65cT/
FBL0Md7Z9ggFdYN/vLw+BGRnUsD94Y+bzAGXKl35KjYwMUWTAwtDp2s8O550tOYYQxs6XIa6IMNk
C/Yp+aKYtgH8gR+kgUKpYkT+Q49RBTb7nY/wd2xDQ40xkZfA7pdJYyKeoWZK1TKZdw1kOQ4G1Nol
PnQws/5HCerjiLt29QIjIDnP7VkyjYSb18cpPNU4x/o4i+fpgVd7a83tqw5S/8KxEQ1VaQatkoRa
wn96WeVenALS3Vbn7R5H6s8IfZbLjvH3XUNu3t5WAKorqQfQczH+ZGb17YkX5AIBKUzieRYTksk7
3L59WI9oa4wdIAR3MQoGd0k/WMh9D9GR82te12azhgXRckJkixxaSDsmpRjq73+p7lyIndrArWEH
31iSm8Gj2l71SZqH68hA9/N73wVIRInyk8gQH+WKuUK7MkwryJoVMnJW3jOy4eRwWVLXzr02Eky8
WeYpBvQfgvD3YK5KfvFSeHxt/i+cM/w6+URUPLwmGIILBhgiZ3hUkJTM/HTqs/zVgFn9NbpBgQmu
uWdWyQlQx7G9Z7PNwcSMcqS8BSKg6/v6BBhvhE0PFUSqfUSdaO14VhGLLKlb8kxxYC64xp1uoHxg
rqxEAwITQjvmh5BHdfKQC9To9R3TqxS+3Pg7b6ODaWCxYyh3xBjlXFxvbvlwdgHzdpUkGil3b+DB
hyq+VIFnQgVdLJ6L+xb3cLGHYuwMH7j9VreTK5w9yJfobSc1k84cNnQFZPE/WNBDckjSa9Ki5R4K
QPmc0X3mAuL5gT1ykmmeGd6Hbp7ecLumz8qgBnCIvmr/5iM3jOHNpCKU/wzH+aa/yF1DypLbIR2D
6VYO84KEZkmOyJTd6RlNSH639GrpAfodg/d7fzzHUTrl1xCpRW2eajmlOGZrYP6Ca5ULTmbyxCXZ
EeWY8DDe7RT29jwk1bCjnCBPJRLM82r+O/DafJbBisPlexdeujvI2tor5NyRclaULuA0K3EdG9fK
7iiSIQD1yyunB1K3yiW56kNPst7Eo5YDFO44vkfcgvzXsDjl9G9NsvCVsowm/LfsNwy3NeChqKhA
EHkuv6bVLY6IBGFT9t4eVr8BDMfgCTgd8Exkou6OmKl2hvn/c4zqdgPMxqLtW327OKDFOsALCevf
/3FTKJg9zzNMON4Bd3qn3iYLM3yxF/r1BQJxVc8bSN4HtJOzwcWVvENda6xXsibHdC8ko+4H1Q0y
yXXnQocYF+HD8sCK6LhJzi4nfmL1H8h1yzC+f0B++m2dU1+DNIrn1VA9rG0S629Lw53/gh36t5T4
ndWytzW4mHccJdX6A8+hciZOKmsmps/PCdDGrUD9dZH1XoDHMkT7J2LhmBADqH8xTZAoMipDi82y
kFm3O6bvQ2L7UYbwKvVtYcOJRBOiWbgNvgu/pjLrtWz05XChJ4MpN1TNoy2n9TPCNjgchs5Bcbc0
6uOr8fzQ2BxKDDcLhKsR7LvLyJh5qmi4l6NHDW2jx4YbqGDMr/bk5kksUEDnJk5eUrvZcZMde1eR
lLFtr4u73ouC2RJL/1I/jYihhCeVWEDc0WPcOZ1BVwxB4Q9+bPp+waZR0NBYAqPmVPyfIBxaVZyf
6Zm7fbvJrD5SqsQsj+ScStgM80w18mWOplH6wX8c4sxyHItQFrjd5koLdqJdaXiPp99wlXNk77VV
IVh7kfHbN/CiZDSFU0juw1Z/RU5l0uEFcPcWaROwd3kDFqoeU8IJ9uMyCA9mfIhe5MihYac0gdnm
2lXOe3fEXHlO141PwCQ3kchrQjxgx3EKJOR7/k+P/8CcL6oNnzMdywzZ4ah7S5iyD6gEFQ2nCnH2
vn9AjK+sPichFJgbfy94Ax8dP4zmYtZF8u7T1SKcnCfBH5wddEGs5qCHUjodhQybfsIhWZJNgXZD
Hu1xcogBC6AovOuekzpf+zP9bkEcV1xOBo5EqcnDaTU/Q07ceIm+hXjfgb2bk0CY0LoOHqHpMiym
i1yLDpAje2qGkvn3mhCcYY0B3Rnd+gWax16wVGYNi+lhovBqSSzlMaduZWLQJUsQdrB88LaYGop2
2zOffpJC7Xd9wBPAGle1RoR0STAOV/1fs2O1+hgdeub6uHU/sEvCGC1q0jTY6Ao7a0BYyvAzoBcg
7U+idRTt1YOwVuGDvNwQcZ3YVEhMqOQC6YpVtevm9+J3bQQquNZqi1YMiRPtCq4PdjXdaSrjjd4q
kqigFwi5FflMA6XTqn2Vp6iuKwsW3OzsefY/VCNpnd65rJNkT2QEwadT+G+gidswbfGNDc72MRee
kRWfwhh6tSp9krRXRKvGJ3Gl3KaNMju8gHEpJ5QDmWqV773MDAiOiNvhAbIyRwpXI6kSKZrloBdy
3/AIbL6+ea1pB9G4pI81E4bRlsF/66VzCsk4VUBxvaBqdhYkmg/XAp725d49X2lFFD6LdMOmBPyx
A3vctr5X81eebMW2H5qi6m560JJx/cOJ1soboPyPg3RhrK47fLAGZnlW22yvhT3pENZbxpVyQkoN
pdjV3S2DqEobbWV/MAOHj3RezkitlXYutFvomTdZ6suu8xR7Z/5yKmS9a7PerGDCg83q/zA+CbFt
Kw+zycMDlO7c6iT0RPAasxRWWUme3mBaXIGWjveHquPZZW9Z9VgTn6Tu64bt4YYV4DoCtdyLBsEC
tat9e+lFZ4z9PWm8SAOar4A3oQBU7TIo2IQv1ww2EvqVnsqi+GsfFIilTw7guabipzVGDO48Z+6Y
UHn97sYi8Dc/Gq5Qqg9QbkFHf8ZCB6bdbI+FQQ9TDciKg5sZJLJHjBSidl8npTuiOCmI++IIeOby
a/2YBBUBcUZzj6/GgJ5CIXTyv4o0SDWtiwr3+oKmedSfx96Dp14n8MakAFuJIXSdFEAB7dTpUOyb
cW3tElM4oek3ffdR7RF7ZU55G3hzUoeczpDFtBiR+PHmriGFUjUzxvjICX71a+KLd9teF6/0sn8w
jdflN6NKzV7UA6tWG3E1JNYR2dCsQ8tcqzyBYmR1MoQfRWnqF+QyWwQY71M5RkPxUgO5XZcqkbYt
UBc8aabtXOuupVGJvuuldDy874oV6bmDKAhQhQbgBqxX5kkTOtOZRgG1tdzM2l5zTrketWSPboRk
7zUzoV+STuTCodlWqa4JL6QtUpkJl94RDM/RULUwsCAIiPsESJlTVk2oCKScCSWjv41MaPRWlx8z
HtdnLssBFIjRAZNHBWP073jSPX3F2FIkrvrIBDyYrqbMFPAOOcYYRIZxo2zFF7erU7A9dDHXG6mH
ESHyxerAkY0hyoReB1JB1FnFkCcWHfqXDYdp0LDDy8wWzWJmFfJqpuq475houEvfbeHi54slyH2i
haRKVz74jcAUdgR5he9ina7oGEh8Z8ypvTodH+ozxdAUx7/Tw9ubhnVpwH7gl2pnRcc1NJgXwfek
AQwiMPg0Tm087Ah7k/00XqzKY6Vzw7u+O17myxbQ6zHA0SYQeFZx7D/5LhzWPRt8Hm/D+nRfgEpD
Svvf5hAhn7YDQK2YFHEkFeXTxGXXdV/QBbRuTeVZgAvkHr8l3rECeovBvFq0T2SV2MX/xs4KmYNa
pEpsFygbNH2A+jX5A9c0zwnz0lYnD1GGZpu+ROLK00vBIA8TdA4dL3CBMfDyw6pw1Jm801QMRgys
/+KgdmWzrg38L+rz25vaBeDTFSq3ZhYToXJh2D/s5w12j6+QXHlnnGmTIIQu6afxLMr0WCeOSkbt
nYDXrMDhzAjW3X3voxsqqo8Po0jIE2I5kAoeZU8wE8QjHj0NaktTrvvvsP1gJa8nqplcoYaSQ2S/
8+b6lJvibsHmoL/MyTJd25kjmLJ6poDSoHlA1uv8eoSoce5MrsLGMmGe5XL9pCA6KB8tHKZWBSCF
B2eHpCxEH7ba5vcZnIYSAzax3KRkmvZfEMoH0DRUih6jmtSYkGhlNRB6TG5rvNXCv3diXoIaOjK1
kp/KOAN3GSbkqN0Zt769fTL9a2igy9Djwjl6KivQ3mvADt5GAtsM8XOrl+xQT21k0Rt29vLjJk/L
mQ8jDLT9Jn+THBeH4mGCkV89I2ZvlaG+m1Sme+CZJs1Der6dfQAIHN8hf1uNcVOjm6yF9CcZZXNq
vnN/jYqjT8RhS7JBHF6n/0Litc/fqUB1wCh7uN21iviEqpmpVXBHSXOhydADTrB5Fu5suP+zEHI7
0vyYOgMu35DqnrzsrYqVJQrm61z0Bff6obTi+yj1reBSc6lT2pMze16158uNtkcfCzB/MV3YlBO/
lrvs4NvMGE4ZmyuEHNcRCSpNwRNfhcvaMCjZtKCXszbR52u2MAgmHxCrpJa1zaLRekBfimyXGOw8
LoFtHA7fVUvQyuh/bRgshR5A184pJN8X5/G5TDY76HbGk4IbmVNIyPvTJu3QQ63srB1Y2/S33Bwz
JTtxRa9lFneQ1h6JjOTutc0VmtnMEN3/xBzBxdSAVxdhd/tcy7eqGSYDSMlQunbuV1hUH0dzgLg0
qkgCNeTA07FDV6rOhmkjD4Fld9wIp3hu/l0kpCvk4pntaNueEvJ7Zq5ycQNQaVREgQ+GCd/Bgb6X
TBjaaFG/UL5mjFDcv6ddPpc9AnTvTsl5DrpN9z1AnDkzn25ptiGCs1V1PnmoZ+CIEYnJwVfhh2m5
OlOxf01FWerFPkdB3zF3W70TTto4yEzTmPX+N+hX6qja7g3Bl7riah5F6mWq1fcSbyEDwwyYGz8B
pk3iOEtU2PIsFrkHHSJBmgMcyJPzvySmv+mwjKC1YrwznleX6Yl/OsAG7JQ44XPYPyFxLSDqQOzo
3qLjXiW723biET2lkZQHtBBTbmdC2BVAsh7Q4FJC8aAlfthHrdDZFgr8Db+Hqt0+3uJgrUML/mtA
X3zBC4MReee2GB5U8cQ3dyJR/7900Z5dbp1YXPXZ0aEMxz7YeEvCVgmc94y6Dw74GVM3Ww8jD6JH
IqyGuihb7qltBSjri3PDPvs5pMSTDNJGY/3G7dxrKIjoZ5yq46fHRFcfXbKaKUIrinn48Ig3VFk0
+NMvwK2a85Gn5WHWb97xF1AoAtKdO/h9UA2fOPfw0GnD7gquXM5kpGtyionOqi7K23JZiT5PSxCU
czwyfAmLy9BYggQbVaT0+HXZd1IFtHEQlnmiewy8c4os+SxM1Wh+pcD7riFfi1DBimo05ZtxOmZI
3vSoTN35kO15XjrbD72MDiSRkVk0V38SN0JyDvVVxmEGrVg33G9C9dhXyrL6xShGBO4mm9DHO1eB
I8d/bT2L+2A0KbKi39dieYKEJFgSjooSB1VaRu1DSwhY9/acbWrCsnJQNSbGtk3toLQEnUoa/Mz1
HHe1ZEofAGz2NsNX/JO0iMpTADkoJ2+P2znSkEzqPQYUvXPBR5+CVu8pwUNQTPUlKkjBGALY1eiu
TSDqHJ6bbL65j/+gd0ph/B06F+sH4vR8QKb8wRNWbXBHN1XM58/Oq/Xhix70uYoOhpLAzVRptyER
jbTKLURDkUxykO2BqMOjKoApGeC6OKSXB2f4f1Tz+Smmp5+zcyi573l+NN9qcx3oAPIOXipdYGBB
EK1ACrHMFMmyQDyWzWTQkDaIo2P2yzg8EP1FMPlLUQWPCp9dB3Y3bmDqP4wc2LY6MfZTLKgZ3loQ
UyHWrDcWRGE3SbeXYMRsW/pS9peAEYMFwARXXzXbmiUHjuIu42FkV6k+SGqOwTqsCCtik+gUBJ1a
uTAV0jQ8qsFwYFnrrmWpSorF/y0h1cg11EKHSlef7e30MtebTe2W0bHhMtKUCLjeGqaZuAuOJfP4
11mOGxI51mpGsZxd+dffXRsUfJq9TAQ9e41YcDnM9hASjx0S+ahKhllhJOCQT3//QQ7pmeZrAUNd
lUwK4aQIGXA8cvHJM8Jsl9MlJTUqphVt3BCuFkZqMoVh1sTZrkcr9IwYZM0DW0365W8KNTJpxEYt
IHA0VegMbPNklL5aRGDagtMVbbzR2xE/xq1XpyYMr61liZ9Tununwfo1FlqUb3tfylCIqssK/OPi
Q6LJiLcLyudIrwbgYpR9cR9i8KUXiQ9C+KTVqsdqdiYQw79c9GZ2U6F3sRDq68WuDtqtThs89MK8
YlxMc1gapYzI9drTZyE4ZG6H8bFqdszWhlZBufwo0paoeaW/WUBAPzAewPQi/28JgxOjniyXP+qc
FANeiU5m6IFiXTXDWCFCqJlXYiKQ/DV1pqjyxYweg4MaVk31i1BiIFuf84/wmmjqBUEhxJu0K/r6
RFsOKjXLma+YaYzabhYoJHKGdGQ8y9Fq519TeZKcII9LX14hq1A1keUT/JjWzejLkkOtBAmTgAR2
nPAj+jAmxZX46ks1pJnEaOgiSBMeOKOX+l5QQdekhmLhdi2lR55gdtHko4Uiy5zRpJ3oV7PLQzUt
jhq+5tmeie9APkKcU6E8E1jrdKfJe3hTLOpNz02QHTv0fCu5B6FMt/JrjOQkxiCk2fLehmUsQxoN
suEL93xf5wd+wSsNRKfOFA5nRtyefoQcl7+Ed30Q0o1XtoDjaMWfc/CxMSLhPTbev7fGwXrcLy+Z
y72LQY2Rl1y/1NSdQIeHFBCsvjYlSvEbiMFzFYgetzM8mCiKOT3du+eAqoE9KaIx0/hDmAOdh2zR
dLDvfDXdZIshaNYyo9gvfBMP3gfvfhAwzaJCFf25lRaV4cY8s45A7pG/5Z10uTtovkYT8eG0Iesh
n1nzZUGG4KS50/EI17g955JBJvB+ckYps1CGLvxZPPhSo8QFbGvwQMRSi36aiDE6794CxikJWGle
QLa11jBYjfKFZ0Zc4Ax6T4509sXo6J7LaEQBvtqtYtWjWwxJpLqur0YUM1KWVBxSnIgWHJu68K6J
1M5/E4dcME9LWqwhCmCf/xqGsOC6D+as12ClAxUj5Bv/WKFiGCWd1zeZkw7jfys4R4OANJzYaCw1
+CHrdeaiWXfuRAK3R+nUiN41y+b+wMXVCcV2j4/tnqukThSxvaAD68orRnF5rD8dAL28WRhWCRD4
njJ82jmF+w9gQFUDrpDma3kHGthvWbqEXXl69di00VKp17P8p55z42DvWk0V+3fNEHYxNoqM+Qdv
73WIoKCCtq2pDbw6EzjNMrh/Tvaz2THrg8H2xR6ZBXLGt9CgNqvfD17dk8JaEt7tuWoj7+PZapqL
CXmLVXqpFJ7e2XYZA1iIhPj3nwjMUuS7Fue+gzQEW3mHlYqWxvixuN0w8PF2iLz69KmGkIDv1nZa
bsIqt3l3tcjiIh23f3j4O9gvzZAVfILjC84ecPbWMdtXMb/M3vQ/zpzEi+rR09hjNChZqCwKimJ6
2xrbHG/C1d0eF5533q7HNL1eYW/5vIeeY1r87G4uCzFz1UWUmawyEETUaxxP61GVXt3V1B5+xzj+
ZWZoE3V8mh8bVe+qWjLy6ToE19hi2/Aqfq9efbwrl0lS9whurjOV+HJg9zOS2qtawuL5rrh+/lMB
1tP3v4k9s/Tde67CxIj56Ulb9UUojzuVhh1Yyi4Tkgju5t2T3CgucYZlL7ZDKLs06vlKaPhLjg1C
prng5CAegoidxj4MnGEFvYxQpXT9K8nM00aUTbceaIuzhyrKoRnXBTqja8+zfQ8e49sS819X8At/
2FsFoVyP6Hd+lk61kFq/kkCZV9gqeujCVsrjGXon6hmaE67y5zAkQViOc1qTRXSBpWf/+szRcpRs
LvOA5RSyABjqITC/og7sygretSs8wWk2NPne1GZ8yocGY8ldWzAIJZxYrSW5Ca4FYfP57Tfz1tI/
7HS4AhnNXZPWjM4xgpEfvoz2B2EgK4mIOeJWzTcpeWxSsUQdgGqJbyhKU5yOHUKH5GhprYopxEuU
XdyMYjLZongQr8yJMmruRBJYsn27zgza99VGXk0oka5kKFyumDF4obtqHT66Ym9KixxLYjNdUNe9
d7JSuTIODWDe8saXV/355tnzDbGHnZDlpWkZ6lZNLM5+BIH/caVv0HjVNP4Ae3sRSqJXswDeLLWu
woIR/tyajns49MHHDUesMhRBCbtA83P7kmzFNJ7mgsvtHg6tgL1lRJaT3wyaJ12c8YR7MPAXlV2G
BBd3ASTyrx7lFJ2821iyotIncMn7qQlun3xAoWXiTlLDEQzii3QNgkjGm2m0zN2ILd6j67euKBR0
jEP/qWSj9eOtmEn9R6kZC7OdYmboaTNEEz22z975WpXgn2yHCiAgBwfL1dZkx5h9NDR14O2TKgly
tcK8gn+9KDv517PqjOMXrCg3iNTnLe+23yhEJQEZ2vwjlfJ5yieY7POP1hbiD4OXTtSK+TCers+v
Q35eFXYUAa4eNo0o9qikjKfJwnEpVfDF0y2UuW3fT83ri+zGJ+NxcjxOUexz7e2N9bhPMe3rdlZV
ge6D2blKU+nVVW6hdhfH+MvKZpXfDMavxBY/vP7PCwg8tsSVp6pwktL7mSoc+j1QPa9i7yaaX7XB
wNqRpjanoE49UZxql5fnzRUyuPyolmiaPv0CkU0KeHTwoM8jahf0dVfLikRqAk5SLAuiO/knUJV2
J5t5FDWXfBeHqgwDvYKns/eWubu1eGdDKx/DWFma+GU9xWpj5Qv2xql9dt6aJf6kwd3o8+wW0lld
9L9ZMj949ONsrh3FoUXWAwjYAZmSrbJooqNK5kknQKyA+XHkxlAHksCvDdgk+ObjtUmpKGBJYdlr
i9GWpIpz1DGwHxGZOceCl7Jl94HupvXq5uMiIzpp1ibgleAm8Cluj2OHrgx9GweBxQ2SudMVvuEX
dSJpQKVgGy2cNk9pEAdwUItcvxWzaXeGG55gTmx12cDZuvlAOyGwlqR9xfQwp/N2m7o/mHTIC09c
45hKVd/pCw8DORoViag0tSrg+YbLYYcXBwknWyWk934FR/qOLZibgScVhXOJKdLX4DxeTo5CpPQq
iGHCQTuJF56Mt1lBCU7dtvWUqTpTBz6k9YgrfNDQ9S8VEzAoIQF5X9OO+vObuB8Z8VFAojGl6ggp
3BkScZRZ01G2iQ0hQnrqswzsuAavsy1GCFxuQYXr81wLSTCB1FLTLbcAJIN9fzt4my8sS9Ck4mS2
NXs3mL+ZmWzHF1EfHcwfp/a41iVKCyMPJcpm3UCgIqzClIqz2Uipd3hyIbCLEftsX0hWWzdgkLT8
FZR6bvB3gLh7PR2FU7N1p2XrCd2b/wSH0NIDGOhsMedMdJ3c2ncrNu53xLb2D1eiak2nkforQFIp
BTaXyggFbwIIAWIWHp0v7KJfQXmqEh3JEfueVSmICLoWTiFKkH+9Wn1sc1R/FlvAE5DXCd1iC4CQ
JeSwoGY47o9MDPQjClNGsn4bpOJiwzQwqgq8Kv4YPP5IgFs69ZlySHN1mn7Ae5X9mOq4KFWuvKjV
E9Dg6754NNo9akzIKFtsXeMMjvgDVm4sJMSsaO9rCjAY2T+NRqJjhP9ZGCdU9L9EgL0uJYF8eg9i
PpYlezAcjXB4PG1N17djNamv+wIqyQmRUSdOxowBM9Sf0NFNdMYGdVsy711FhsOeNZRYB62rkDP8
jEVnb2/ILsIiQK7pwO+316RRQuyJunbdzCLrv1cNPLjxgVmiikAqLI+PytG2farztVK/eb9lJS6w
s6iqE9SgU/YlgsiPuqWTEDx8z8AJnwrXcWy/oz+qTsJHqOFkWRwX/OI/OgAOPzKw9R4VOujPSFEt
f0XKGHh7dVURnNqeZdaylQz4DUAcmVX2rhLhdYYBrHzdBwKWLkqB8yZbuePx9J2AQfrOdHCb+eil
5gr7VymjgxzN4+FWqVB+XWkJAhSUag38LAOEk1+Bb7LpeGHk+wwTzQ7apeeK9CDXqmcSfPEOpQ1U
GU7cZF4baBNkFwwracrelGC4qKGBNYroyP5Au7RwsEvoBV3oEBFfyalVgjF46mtRULUGPqmgC+1X
Oxu/Iu/FzFserv9Fws7rsWJpD2Qt/5iv6W7xmNrNVZZXG06YIn+cJc6Yzcz36D2vpajOJ49xOZ2k
jmGkXU33nifNaW0hcYsU3hLFJ8CbBFEYsndFZB1HGPAnbryek3bw8cExIfEFxc8Y49AiVr4v8VOf
ZL3/qLwJYX9q8CB/KY5uUC1zm7qLaSBzkzZ4vCqIBaJM6vAHi05g8GfAKXcLfDPKIR2EOVpMV9jB
tRzkejlErdq0yVNj1nHgApJh7ojf1XOQW44Uw44xjkieDPLkO3m5X4q8ScamzCPfk1rKUHL8+j69
5AfwVPSZC4rgFrMLZ6g8Rtc8vWvIkv0+j+5D60eHzJQH6/bu2rFgrwT6TjTva/1D21GWweEkcFCZ
ZolzKtE1PXgnNPLZlgPXoYOdyXwhTQOyvOmJ+wlxYPxtQztO6iHCL+dFiMTml9r1ietIcNYKFf/H
72KzeI7J2R72WDdzffuqFssquLM5nz1ZMSv9Yhp+T5x6rqcUGD9KpubD/daqCPSn5fHQS2jWmzdU
ifX8VDZMUWda1t85b998nVXA4GJ7Sq9X4UyMooCDia7vf6luTYsvGpA5UAEs0+OTJxqTggEQoUTk
LXpTk1zkhz09zS8+V/mfSGbMZ3X6++3+C2vu5jTDQHALbw6MULV2ZFUDeUrNJllYbgjuoyBWswi5
ewn4MCtFaIYsgL0o8zh9wS+C88E0A6ksJHfpbRY3zm94bN0Q5Ld/soQP2TQ2kwOaIzRoPVUpN0Sr
6gs4gTNpmOCjlwpBjGgGUqloi5/TrEVNcx0Np+Wtwatqj/lsnhNjCR0hGWQ/5T3782uBxfWJLqVv
XuRcH4/wDpUmjJqtQfyDqBjz4jtmuTOsE2HSQPgKBO56onsnrIM+hiSYvk+QGN+Y5BJieUUIpohx
zC2Y5nwJthZINwOWvvURWnxzYrJ/jcAr3RjvOoU1guvMgnY4TX5AfMXvdj61lj64woAfdZoKlyj4
cnKa8WgcmAEjFqaKkIoaVy6E5eIuXcCXZVzN6O29gDZebtmcefZEeaMZgMApzGzqQ3GVLQ8ZV4fL
Be5wAgg+hMTe/KunMlXVK4XbSSQLry1Xplyio7WIQJXRImBEGmwvAdw+zl2liDOmISV2MbDH9lST
17YipGyHLhuSJgFPDeJOYWIfxVvQAYh+JAd/pBGdF+PH1tSype6VOtLlCQ8zJaA4Z2XzJDzK6BOl
3eb1xdOISTDNM8Ym4+aglPaFlAml6+6TDBYnQGs6mVDyQ/fJzBHstmZXxL+Sh8W4MCIvqYyVO+Ps
2dsfmidy3tvuHoBSZk/quJMPeXQpZvQPowzGkp8f+VOe89ssnLaKTBngwrQfKeO7Wx4muGFNBeqj
2GyEwjwBBCaR+DsmsjDvT/pzYkDFhPnp6A2JAzYZgLlbtiw0MpNnsy9F0BPPeqKyly3goxEjOLlV
a5RQq8DBNxxLtKJDJX0E68mLS7M8fsi4PeMCF/sJQDKEiqwvbfZ8/YmtXz/mvI+SFUDYY6UeTAVO
SgxwN6c3oxOg4Yq++3EgpgZnP0wmOTi4UjzjE8Z5Ejz6Ea/g0lAiITGHfmgg17Oa0na3CLoeHc9+
y4HaNLm5nHF79nlBKVaTyRgpOXOEm25DzqxT9Oi86/eBF2pIMXaVad3uobRvLZE1wVIiWrd9Uhd3
VSkl1PAN26vb+hoBlHIgW8ruB0dmm1hz/fXiy0gyDMnrdnSjrWngRRdMORNnm3m9OKKzO1/YTW/I
UZ+kwbcpkiAlK7/IZXjulsja3tUQcotTuRXjS1yWT+BKzjWW/EUtOEp9b4p2VgDmv5DhpsC37CLF
iq+0cuXUhp2+MipgHBA75pGB2KG/FUCBO5CzD3rOm9OGFGg/SceA+QMAqu6vgUiMRlKHjoqTkvB8
EctPrK9p0iRPqjgG/t8i71EUbtV2dZQfJ3EvcMH5W19sDx+8syvDuzCkLj4SatSrhCJXJ5CBLVLi
qatxrw9jow5l7HCCDwKudQD4IUIffjSdGh4hMG3/ix2FAP7bMwzNLWAPkpq2dAcrLsUD/I8bzy8N
krm9vSXnrvkVB4I6/5cdXeLRzyhuiniTTBV/IvOEIPewImswEeR/f31UOUjSRdKYlnRxNJZ7ytFv
X4K0/fjtin290Wr0LFVslFYdxOMnRS7TTi/R8oVLvSuC8lE1N7eiDdc0OvxM5UC6Fr9iQfh/XPaF
zIrpvLswQMeQaJ47iCOKkdTbsW6PpEdHOjwiflTPq2yyiUrDtox9MpY75HvWVy+OVzl++sdMlKAt
croqkRwbP3dJtYbemZ9TikgUwXzf0MutNgOY3oRUVkNrJLMvQ8NN/DxEVkAohDS41p0iZuJxK8cU
Y07c4VdgS29/ZQiyWsh3xWjkgnRsGdMNuEdUPNqaYT5UtD2HCEE6TX0/5sWYdxTdZRbE2bTApgCT
Lj6wWkCjeCCB8W82HRqAy3GMWprYtq6E9rliVGJa9oTCWt4Guveyo5QX6Ymb+/rH+2N6EUSUTP2P
yacJ0mGKzwdG8PnqfJphrbO4pmWTYOjmpHAFG2ahuEZmqWp9xNu5y6LaK8gdTX5lnfKz5icoJ2/z
bQ807FUV9rNMLt+znBz2ZrSixzc7Yf3v7bsDhbEcjp2tfz4pzTqaajAdJ4J0rkEey0p/ndHPN2qC
OWAyF5OLsfBs0TMXw+hPB1ippH69nXsAx8NWbhuXae2gZbPEU1rUFXKRTAScdd34+ByIPz7V2YiI
ZQU3+Vg9YuhWUWPh6MKUIbJeBXWKNfiZJM1HtI/MvEym33ftS0yjcKD20BdhbQv6GVTQClHNLkx0
KoT7QaBNJhg9YzIWWxKpixg9AyYWfwzKb3uFxYRnrjvA7IKQs9eInFpimsN1ierj6JE2l6nuLHlk
rfnxdT6VxdocinHPcHodqWEOXFcAIyAc8rw1NidqjvYBUJ4qGUjZLz4hNy1mVN1XMVkFCRnobEGu
O9N5INbp7J2VOFjZiXVvSd5syVonomb50UicZL3wJUWyKerLL5QdzQR6hksaXyG+ZxAqkIzp1TVO
R5bDw8LU2DURGplz8JNZvA5GCsRaVhFiVUs0e70NAT0hTJGAkWIBUXRFTgxIfftH/Yw5rALTzIfv
ZwLoxeF8DJZQpZlCXIZXnUG8Gm8FzLzGK292P5XRvq4sLmTWdtq21N+HA9cqOfTldmNb78l2Vfs7
jmaDF9UWxXMzrKshVS8zcxnKkDwZeoQhxa0y+u/668hf6/IZMAUqTb1QYENPAIqPh/sORUS4DB4f
CAOt47aSMBwDiWYwXB26mxQyUtColPIsJik148ikd1qmZhKmdnaohB5rM2vNpUcypMhcYqnW3Tuk
p7hnVfXEZYxdcFzdinWdKs7VJAUuzyJ4mDG6m+cG0ALU4s11det4oFegJD5UOB4OQT7MCtbgqlof
TTYDEaSxWBO5jfbH7aREfGGCAEUpe6whPZXc7BB70lsoevWKXP9p+sAP7Mk7N1c+67Cn7lMZr9nJ
Z0JYrjdULFnExvlIoroJ8JdPB4V3m5g+9yQGT+8uZJ6TH5thrYygjvQhu9Bmw4RCuxDB55B3g1bI
Fsbxv11A3ex2fFmKaf+WJkydHuh3ZEjZneSxtbXs8jzavXiiZnkoYNG9Z94/OY3yxJTYw5wXt5Dw
1GjQRfyx4zLhSt7H5F2xMl4agbEUgW/AYIlTbs3vFw1d6idf6cwb5QubcnluGT2De+Qj95bR5yHj
xAz6xYAOXrtj/mjeSFAzip8HUt7A8CuLGpgggOXen50bRbBL1KkQXvVCju41+c5UelKMwPYO96RP
byy1QcnGAIGO6P4WtDQ1JL1AOm4b1I+0RTRnHw8Yb/XbwQJ5ncIeO24I8SY3BymhVasVBj3hziak
/2fRG2XIi72ujkUMh919kyATudV1RxtPWl8AJ1Ea4uC8qwdeSJHWUJSuhQA8AzJFqIcV4NDnPNs0
9oRZUgrNC05MvDJoHn3043m1Xr6oKHcs/W+w5GtKJSojp6d8zoQUT68p+VUWUuWqHSKT8fb9Rz1m
QfmFJzDIE0haXll+fJdd1MP3WQqERMjVKeTYKkm4TUAHgN2geZhO29Q0PrhH1nenH+/0Cv7JB/Kh
et343wddR2LoJ1D+mSH5VGESzOWCj1bzkVNcd4p9mal7/4/4nnGYteGbXVNWY6Kxa/QqDYSDYsw1
zLMdpmH2BACuo/Qnk25DtBBB5KwlM6bGG0bjU/7OvGAZSOO+C4hxqkfdD4a1ijLnNrByM10gJjU4
8KZDH59o/inmPZfoxar7iZmm8tKUrsAufHNrC3C0gZSPKZupjcZkeIAPwssDqBqZW1Ek1KV4+Reh
kQpLcBrOYOelk6fYAxLN2Rjj/IUWzy/sr+l/PlIOvgx0uhipcCpYV1KCqiV84XKiM99hTn+bJR3V
k/wbL5sB4SsFXvBf9XVLnvTId2PT46tcCxp0NTAL/NBnNHnmUn4uOzyDAAyi3Tq6lrruQW2htjut
0HTuLGGm7Su0FI1s8ekYbLH5QA5dBlIWTzbOi65U1KhNWkWA3rwYxS6lVYOy8wU9jEkyUo7Z6vDe
CDiqWfz0nQu5uCbhZpgIrVJb5Fj29VG8a3+TlpeaPahF8Kz7rhcyulszUmFjhRMnFtH4Y9wMP1yK
f1uMlBiPftULDWfdMru+VqhBkpO8yn6V3VxfRR9YiySZODXViY/H0qoD2V/lLkttIm0J69jtbiGT
PMrDa0Wb+9+gMLlNYqA1qte3hlAVlvTBatiJsK1P11DNeNSDGMQDRuqkQ/od69LFo6djep/avYze
oWebPoZrPGtBjcA0tLkROk1VhUTZX8FBrJQ52HJmvyYg5gMBIwy+MZbspPYOjILOjM+S+cPhwCrc
DGFCTiczI50VgogKa7ZuwZnDQn8B31csBravnuA2Iw12J5LQ76TWToiHla7Jtp0BsKfZjGx+psLb
KhBmhgMCy5t3MGSfXe/2JeTAmsKDytc2KpJrFWMx9jmyh/lDEt1Szwb0POmtSV0Sffx8I521WVRf
W6vP9IvkkfNI5rUDvL+ovF6/9TiNKsBqA5GYKG4MwRXMbCeSTmVZUXUOhjkOrWbaaIAwygVUPRrq
OjCf253oQSj4xePqfrKaQN4Kvijmp1VdlGQp09syHqfcr6Br/o4jJqXzzEZL4iGAw9rZN463lz2Q
NDmMHtqsaJJ30Pucu+NjZXEz2KQHRaO3Ct21ffPEVdIha7sBM4st4PWPb2dLeX2J5uHB7SdYEBYZ
j/N/awAf0jmJ0MoLI0DO0oLEQdx9kdlQ4yjplvIR/hnairXoLEoU7wRGbKdaZBH6FWoTXybWEopN
M4XVBty5vye7k4tCCE59iCCMFLZn1bwupbwVitAJv/djiEOqk/+cAa1hMdlDqchk5G5/1LA2wU+x
ihV6uj7S0Ioi5ucGoen0CW0krGZVjbxCE7hl3a1y55wE++GxPMcUsLNYdaZZyjbEWkO38O3OShEH
1EXkYHuUdM/LvuATwLyBwcEpQ8WMvk9ooWBv9oXfMMP4CEFrGGrfWzU+tU+8f7SxNcYP/EPFuhdU
jJF/3xthIugfAU/to4ZCsKgr+XHXbf2HE7SvOzM5tDP2KLrm1ibOGyC2A/9oY7pl3DTkq9B2KWYS
g/l3WZR6V+06OsBRn/BPDPVx1NM+EDemW2u00r+OJwdRjR1OZdzUVeSIwQM9GTZt51iNyRyyTs48
RZbGBYzR4Udg2E0Vgvnf/4bu7I0prZSpomUfCogtYYQo/VE7kdRLQ2hyjR327HKLJPOfMXoRsFQ8
Y4NOiu4NmHLWxsys5+mVexn3AG7mftZM84vlYvVGcctbMoQsi7V+Y1XbQtfHmfuCoakYbImK0oAt
T2EnBmR4d/OzyF0W4rauzuVlNSten18VYtzw1f4zOHz3EJ7fwBmW/BRjzOMQhXD+NlA0+Jv7U4r/
LtKtbaY//esNcJQitrPB8+XxRlRqkGuajwSmpWvnxyQIPiV/9KfEPpH19YEXPbRm0ioWdBLSlLBs
uYlb4scYYW3TBWpYIyWt0JWgIIruyuHoXTsTzQSqIjl8ImrMFrTiHKY6GSt5uJNaHLmG7eK3G/Ph
qji1qNSn/2o6BM1T0RfCP5HRQ+150kz8Ki6hmgSjaSL3w/j5Wmvc4atCl2AOF2bKqCW5XBQYmWdT
1Ld5rpzQIs8yVITpODqHiB6Cf2U5b9nFYryipLpFgvbJUzFjsklxacZHEvDIWrEBLt5cPxMW1Acq
IjSeWWbYphslQZeqHfMKQZdHPbLE4sD36ziScyQmrzZ7enqKuqKluXsH+uYMWTJVVx/pRCzBofLX
k/XHusyzr8OJJqrdcxEUZ8di4SiaTE0fmgstlmKvMOxpUz6Tf1GFnNE90VFxnVYTotemdXNrjb/L
fUiqftvWb9vtQozosbHeFGypLi9eTP8Hb8++4V0/Pawbjy2l+FnA8qowYpTjKZrE54uGsrHNMSXn
WxLTtuoFdnqE+bB/SUA8RE4Hwz1YLwypn/opAkQbDoETU6arALu+2O4eo3s3ZBlf1XL56R3XPpvd
kqtWC56oSrsUUwkNkS8ln1BnLgcdFwBgyU3OMX+rusBW2G8L8Y+yn/OFW7tBjxRhZCmQyOO73jXL
tVXmcvlEySb/Gmq1A9p8qLUc2E9DlWtvvaEoRjkzEUNwDZDQGrAR+QIbOSX2lhQYnv8BIAeon6Bg
ayYsAqM1mgYkhwc25rQIZWoIE9GQYNN9uamN8oNuq+PrkQ9ilEJTZ2hk/qwMfvsGXVaEHHg1piCS
NCSFsg2A8qxxuabxC4y34rDFfPPk8og3Ha3cGBvS7ytpSyIZNuiM36/MWQlE5p1o4qKCqfrw0dCN
aC1tkYzQdPoTPmgitdAyHLDog68SCOf5oB4skQv373CtEdrK+QyTrIf0J86pm5QVijjxt0PvqNCq
k7RfeGGG9AmIg6V8fmrukm3YY60Ya4eJJ3n81Cps1KYV56KnK7BJ6/kNoWTBWCWf+W79V2rj+K4N
vJnRMzmu6Md1WQ76Hes4A+PfhBrmqj4td7pX07Ndwk2aq2JuZ3sCzPeUXc7tz1rc5BrE0PBCzTKK
5Xi7P/ZI3tFsVGs50HjL2Ns2xinLGoQRZPqeDBwVTYqkRFGn4jPxPsgf4xKtsvcgFnlQrZGfiu1n
913RRLF09egWzQW80TM9YD5CbxcLN9jb9+/2DDAZKRtq5gwuvdvfrOGMmP79bLCHGalF1/Y+TmBq
SIs/Tsd2kMFuNqP2fJmbkiW/0z6c/TC82bExnCiHGZ0EPJkRXnqPvskGHmu32ZTpR/4DlD5sm9iG
Emka4gZ7RMiF/zfUPByeocKHARkjo2WR+WKv9tEkJxsg3MuRVKNU06lDpNK/qjBgoUCwKiNAU02t
krbX0fIl4bP+ecoOeYHeYmgLcbX1sTts1/2/OPkgAiaHRvz5ruE5IjVkmJOsqIY5JelqfeIM2ICm
8EK2DzYfIE9KknYM6R11+07WlNVl+ZYj0zWhrQeAzEWeABMoFqE2eXPRjszCfBz0MTHJK5yotB9D
NgKolf8ecYtKozZV5SUTx3EYjbewOvBFQU9qj/PXcZ2bKMLCSbdcKHFHByDAYxDTvcynA4jTxw0q
DfA+zShVje0uTzdtWFMTn3kWLpujWutxxIODyl1U3lkHhEEStRnSB0y+6Udko0E9s8Y2X4SNiOPx
Var+iq1gyiIsDX+PtpZfMeiGzNDnimeXptMyOiZ4R5zxp7qvvOftmP2u6ANQt+h7U41yy4bAjEgb
QXvhokeYuPHi7Lp26LJFY57AYMY8K8SFZUT5IfoMmt5QW0KMvqw3Ku+IW9qMtfFy6DoRALKtz63X
xbr8qgKOZYzD/pyFgReHCvCe0mqwdgYuwgjChdPqC+0HfEkA1FtRsPKUVPp089+QG4T8/S957SYk
h/3S8YXypCnmFqirG82twJtdYCXZTM7aR0QUxefJNtwTJa4gRhCdDLWtraa0pVjtIlCgi7zBXiX3
Tx60FdyMZOhHOH0jz+M5/2W8jrQ4oqeiCcM6Kpai8F6Ty++/kM1kRQtOMxg7aOzCUu2GA+WYvY4r
kAehXiwqB4EA4WqWKXznJpZxpHigmF8xl+gmq0xrE0H8AEMIKdyWSUO/h4gi/c5Gyl3D8lgfd/a0
uytDJPGEcAfhcOs7Y2nk34n1TeUO22HbwuiLN2At6fqd2Ed+Nb6S2kKyvfOR7sQ7u0qSDxj0LIW5
i8z9OfHrvkPyJ6PeA/v5xl00HBsZjk18g+kmQm3QmEfykIy2xoTGWopCE+Fj987W0DMn1cfckLrM
Qjz0TqZmcusYg/4mtC6EXd+fnQmHPxmM0N9Nzj5WodN/1V7lEKpZSsmTwviDZUi0P4SlEcymkQ5q
qMOfyIdoJrZzUcNrX2B5O2inw3n5myhWG3sE1ZDpHdwL7tfLc+HbYuq3r3VtOmMVKnXOw1vCDDa9
6YcLgTGApK1xF994mVcgRLarqgOxDwGu3VoFLI9jdCt+s2zohlWazuCb/eNyGZdGuI5FtnbwD3LN
38RiAklTgNjZtgYyiUiUZGMjwz51OLkAcQ6CKtKfFodM86/Du/n7PpJQL53cJn1agZvWsTzzxbuu
R8/Ca/htO2Hv5TnCugdtGP1DwCMeA6oLhIRt8K1FayI+F4WEk/cot+ujAqxmf1J3ScI/3RJ60UEi
fu+pQZ2e1D/eqvljVoMrJeQ1sH1LTJ2hh9/XqDRTzlbRhJtXkHqUabnae8a0tGqC08GzHFtW92lY
plTCae7V76iamG/qX8ITNNsQqpF9U54bYQ8LNWtK9hwaxf0QhZqF6p0pL8ni0G6kz9njTSKZ1xzz
umdWlqG9pDjBSF7VARExhp4SazaU/K3MfdDracifvrmJK5yRTadDZkP2s0hc3qTWX9vdCptgE+vf
fnvnfLBYKspVoqHGIzlE37fWfmmO937vlnaqNohwhv2P6D5fvz2Gw5Ci6zpke8+/JmnijYDrFC1y
2om/dFeY4kf5XiyCtGpT+HuO7WdV2kNMr1o1LXvMPvn6LMw5kKqKYXiaaAuaniSzC05jK0ZL4c9P
ZASqKKR5ioEz//jaymV9e8pg5GvJ/cFFaIR1hvsG1pzSPFxjJ+/wREs+1gmim+RV3dDnAz5QKoJ2
vl85tJCIUNdK4cFJiuzYm0gtanAtd2tZrnRQxA8+cq/38HZESt2/aKKELvE/PfsnQgy7ZRt+F8e0
+QlwMjuUDmDQvSgSM8Xi2RE2qQCAxbtkLXfEUfKEOXO6MYUqSTbE3CVvlz9P+TKJ+8NV2RbLB/aE
sCElUZnXAvCj9a9DsegFFZgZWQgbU9N/N7WWrMF4GtiAklI5zf+cm308nTTn6oQHw4dC0+XHd2Yp
MrPFrsvzGPtAdi/p6BloEYkz4T5fQlJ4msKHBFQPgrWKOOYnEj7QcV8RrVJ2dc3sInMo1N3pnXbn
6lWQfZzlI2Nxf3xAwhQ2C6Z94p6AEzYZMkj+SxwJlD0C+6HG+szq9bvDZtR5pEFZCkvuelqSWiI3
8qz0IfRSjFK6RDGIv8zxYsU0GUINNwpbGrW9yQnDkd5QC2L4mf/1YxY8LtJPVD92rBAqnGH8Igud
RTubzCzmyru3xT2tKrWx6G/qpyZ0T0YzKopcSobXePwh1DCrnqig3KWPrRj7m7zgOJhPoO7sBhqn
t2GCbhEyyZnQU1tTSWt1VwxYX+XA5rx3/CDDcbESqUyyeGn9VAIy85hu5hxHg8y/+OIwSVyulOVE
gwT+ujM6Yw2RWV1EzFMgXb4yZEc8t9An1vs4Kzjh9ciI91QzO2ESx1QEe44KG0Ga/o/izfQgIa8S
u2nOVU+jDU55bsIZsfje5llWGHma5m9q9B87ifxaLaAmtTf644rG+cu8GPDYcrSFCd8p6j8Tk+Je
bGKp+N7KCBBTxXIOVbJbHHVrLyOIlVxR70fx42VAdeHbq/yyZMQFerMcgkE6hYKpREV64osm7VuX
+ogZEcT0JnQJSIM7cOhJZ1tjAjShedtlOFg51skDNrDjfbhOsYNSy3TPAae38sfLJpZsfOKmd5xK
ajkJyCnLpFO5Y8Tn7IFrnHHoDhWtqv7G4yZ+a5dDcmLv26fwtBFmmcr8MUqN38yCuXNOUa3eDqzd
kDTz9qCDB2o12KTGCgwtfaqeZIz5cqipCyNh/aCAofKoGSFSBGheg2IJNMjZOP8JmYuirUMyg7Oy
LLQBVOBtq8LMd9mvbeKcsYlS7CTuSJ4b6MOieCTmz0VvYxi03SPW7jbyO7i/54ruFyTHS1eHnqge
5Tw8vapzIHCAbaX+o+CcneybKO1mdjIwLYOSNNbksRwBkdb5kDekglfeo98Xn9n2VLFxItFP/li2
zlxdb0vNAQcf7WMgSgypGJJrr2x/WSvTm+xxcDnvo9ufoWL4BrN06K/W19CTid1nxZModraP80a3
dFSDKPnIJNOW+twbAd6McKneZVgx7o8lrgJy+kOJHA35IeL3DLljFZhxrbB8irbsB/45qvt8diCG
97eutFDAV90Gao+3tW1eodXJcUjFh4nL0FyF75kUNzYgVrKebYJoT0TMTDlH0k3wrjncrxR19pVD
Gfd0OKmkaz10MM+PQJw6PtCMnbi6+4sKg3Iwx5THsEdWGNyLE+RnB4SxQsRywc4enQg9wd4Ty/Ln
9XHwVCGGo5wKpbn4D1jrbktduZV219IH2rCpfDBQCrEZxnCopeYJ5cfowrV0AHDjOj9py140B/vW
EZt5KVurXCYfa3kucy4ZQsrd3uL/sanqVNBwE5p0zS9/ltIWqAQIT/WfUOC9NleXXsWfJejKTqwR
aSDNaeUmfio02b+R0OD59liaJtSMRqQmVAj9wAqZmb2LE/mi3NpdZWdew3FblgbPPnX8CQMkL/KE
GPAPAJedVjCvbGlehppmjeoRmtOQjRUznZgwTUxAEkwY1aCUXbGw9DlErsZ5lumqOxIzBZqFMpt1
MptfIDFW8l7iDqL/okwWbL60gILlDgBZTJBRscoE/Rz7khUmFVvlkT6s/1XhcP1V9XhP7483akmx
lRVezUt7IRc0gTRw8IuQPkhZS/dzP9VdQ3YPpVLqPnk1sEts20UQKekUbsobDEO2dbtfya3+lIq4
RuRpT3lBSeiCE6ltQHaG+1qPRb1wRLKM2oExK/xSUtP21yBSZCKKHxAgVLQn0DIJz15ZCgwbrR0s
UAQkmwf/KT2w2ZaFE8n+SLtQpN/qi0nszOLD6Kde5gW1ckVdlbUIqNHAAAZqBigYemHtaaRmttaD
cYChbbWx7U2D423oMmIRCzaP/Nqd2/4o37NeGjbx2C+4ywjnUf0hacNJe92yZ0QfLTzmqarrOBt3
Vzm2PyR1iSTh3pLpqafhbUyazKVfFcutD7uS+b5FCmJ1NeTSR6k+ryREodpIEZdoWufjmvKXuw7m
sg5GqQvPcRNWSYwy04Gbg/RGoAjzGHRcEvbWhJvvzaRsRGWPJtQc2XGYiXDFmgBsc5cYTsaq+ioF
5UlVgTiSYSbR27IE+3QzN0GBgHFW3jUiR32toJhq538ZUNdAaQ5zbojkCRDt3A5toNcEaCLuTD1h
/k6vUT/ppwJChwH+DwwQCc0kHyxI9QqUJ5ladO3bvH/g8n5x1q+0nExHNTW/CEL8euV+UeHBezoh
JLfBGZTc1fYkotfCo1wcPlQBOp41cSeK1H8ZVRad6u8SurM2CSpAi2/jnxzYq+1vxc4k7XICgrd/
aGG3lHLcFJhSIAEjrs0Fz1Ih3Fv3P3G/8XruJwTdVWe+kNFZJxAgNdbUZ28vRf7UuAlrDF69AxKB
EUl/vjPgLFNJzsZPTv8Wj1hroSHJa9paevYpRhi78grYYnq9DIDlK4PafF72H11XXZmv3boUnc8+
4G0vd3lwph9Qezvq3KaAVsidEYf3rVaByEqqNglQmRZlhy/Qt1Xe2ZPorEm0FBG2y6fa2vQJ8qSj
sKV9oQNZ/EDI/0TpObyW+hBPZmAI4vaKQmYc3XZvv4cMF/6Ok1MHkczEtO7wVPL8e13lvan+fDQ9
ki8Fei3vC44XKnZRS6CacN1ULp88mdKt0Qv+hiev1NyMtrTr3jlGf9/ZbYXyI6ZgZ1plpsjS7PaM
tDXjM/u4QECDurTfvyLJJGPdzXSFLMvL/ZVM8zAdMGsuxP1cGtdGzAAjVcMNGJInKeb1B4xLV2mG
ENyCiih7pdBj01BfFV88OKtTqk29bamQ9CP/eNzE0hedvi0to+8bX9C+C/vkPXciT+AeZaUz2ZSl
TKv6lHxfog9v0VnLuimgD17ywPVr8x6kSv1hW5VN8O0RY6x+DCWbFdbhBxx9s2MVb4Ja5et+ye5P
oD319woPBHWQUQ1EBo7CqRGxmB3ZAwTnNNaqZ+T9t6tQFyX6XzJMmEVTVXNhU5vRsJBC3oXBGo9k
SxwCSaKBdQgOFWoMvxfcQgklVPVzDlTRwORXw/ygfeanhStbwd10AJ4cL4Vgs2yTzCS9USpxwAMI
IoixdT9pUT1IE66henCSxOcsZHClrLklonKRfg+1NqISAJ0PeO5X9uFH88Vptla1yrw8k7zzVxoE
k0oWck88xGwuQm0gK3Zs6viSF97y/5eWmtWWGkWmZCovhi6xXb3g+m0Wgn3WBtMPrDTcxJEyVYQv
laIns9JONw1i91DfFRuARto3Ad5g26OwnEFD9mJU4bmTX/SDF6fGwTRybV8YJlbu8p8i/gsgCr/f
0j9SVPtC7UWkFXGTkNNS1RaX0BjPYDiG5wKzkraVVfNnFLfL+9fApavCIwU3MpG079PJ/HNscpz6
/oZ30kr0gTXjQ+wCad1B9rhCD3A7Bs0quadZqwddh7O4gKoMrpQKb02DGxRKM/knloZETmYM0Fgu
cxdToWaVGC+DJvVZ5Z0EAQvt7Ocuq/hOUUNFpAuauSFI/Z+PSNM5oBdF1Ho0oBLT+A/oVEvuB7dk
RWXfbqM3HMeBO96uDsdDv/A/AcZsHscElIQ5VU2UL8sC7jnwejYixRKr2a/PZmLQiN/4QeSpXX2v
uJIMxxktPCYsqv2Y/yS9dFankwONOK8/nTJBkMEhxfKoihlW8t9ZfxTuYAzQMGdQb2LeSg6qKyzk
iKU2wBe+mBm8AwknG9GADwuC7Brgosu2zrMl1tnM6QvOqxJwIfd8IwfFtdAPuR/cLzeukdJHiOpN
IE6Xr8U/jLLC2IyZUWfMAfa1Jxyiysj4QLlk1AzYCycWsyUYb5/ajcZAPpU8mw/xYXf3W+93LRkZ
54ANc2xOUhR43fHJe9jqjquk2+IctqGl/fH4y3sxLQzQuNQ2BEgw/r2HuvXCSx2Ku/qd2oXVQknb
q/Jdn+VKLtjH5TFskcOUW5+WBQsX56bFPNY49b9aeXFM9W9dMvYfZ7nQrCg9qdemls9LIgswsUu4
UOpv3hH2NFyBrhObkADidasIZPYkaL8yLTgCtv6My9/Gj9UvC0Bj9hkIdNVtpULwyjPSiYVPE2dX
HJzxVcc22ae7tDC+rVQYk5u9jxUgg+SaedJGxIHxZC/zXZCSXv6mnvEk597g3crVdYs7dg8skZXf
4NyLUah9dYWXKtFDgKGJkX398KAg4PRUtbDGw6MpkqwCRzF5iIlhbvCQ3PNpn1tLwbme+wp+Z3nI
K9GjhoC9ctCiUsMaXIbh/56u3O+HtTTskD2mP4iEr48ptLaApupQDQNApyCjr4Zm69gmpw2bnRae
wM1ROA2uvxDkpPI7Sc7hYbO0/BJb7VGLDi2NpvlGjtvV/2kOA+esbgugM1X8Lh7xK1cse+3yOc5w
F+HDjvYtjg7bITFoVsgQ5ydrTX2dYLnoiF49a+MGXHWVFqqhwObUy7MDrd97/w24zqmRS0rtg8zl
TqSAW11HKX6rrHetHN/QFHmtL6BRKPmqxUQeWSfN18BggnvYFIPTCE8yXGHVcElWZa6kgUyy5wHC
cObDL1Wd6sC8CCfISo3ePiZKw7hrNUwKLFZMXDSnkUrWlSnTr2qkT4+yEG0ExFnvO3HjydSFpoIt
Zgdg8c6GSQ119/ilZk4rxnTDjL1Udsem6B52TpJN5mI13mCZq42PZwGiSZ0FNlOsx4eT2O+7sLW9
2HqJll72gO4Il/XOZTLCcZw3MF9n2E9H1Z1vbhvPhT5jowLKhN1AXFLpzpcrMuW4+BC+qIIdgtQ6
K14hOZAgUrW+0gXWCWB0+uoMdfiJQLwUBIn2UmiyO5KboHrVgxL/cGZUCKL+n9cWTY68Xv6iFe6d
Z45gqa1eLEvpFYpgFATJ80hHsplsuOrPziallKpRBQ5auwtQl8Kht96Z36T0hg9gWC1/THt/JHVu
ds7BOc0vux2wPVSTi390qxuMiSaDBQ0H9a3GhwG792LAsZUSg4qqHXFdM998qJLbeROzOpLWsWc2
xN+UsgoqgXcKjZB8sxClrpRhGpYtA7Giax3g0fTRkB76OwLxTKFd19oSZP9LCZ3VJ+usYuU8VZwl
a6pBzWcTOQX/WPdwQL/jWT4wMHPiYSjqVWNjWLyCHyQrCazxpWFsqCianqmkJRbXSBXwN5rWnlT2
81//ybYWE6Rmq9mRJ5yGTmZV9/QDJTho4fDn5U3lK87C8W0oiE6/9FUw5OkxIvYj3eFyt85FpKuF
g0qDjg6mk+HFIz2ADblSi+G5rPJvKCcW/nmpd09ZLrXUrR6d2po75v0IRNLHZMGxZ0LySsy+n1nP
TmHTAu08UgJ3hAdF7yWVLkWiwkKYWaTaEGT/tY5mj90s503TCRtihr+U3s2ublxwT7diGqJ5U8Uk
XOheUPIYi1+8yxjysSsXeXisjOxg3S0iezfrEDx3fBpfmfZGSQ5FfvOimbl6761nZEJixAaPcYdl
mCkA4lHcvFtp0dkABv0DpIScSAB/qPUwR6CFGfvVXdYhB6s4hFS0j+cy1UOjsZRk2riKRVvYgx/y
c5+sv+anL2aY+IZnrVW2PJjbCwzvFftiPlYegOnH4htigL5HaSR5o6mGo22dFx4G/uTdfMTUYXQL
vc90fjrJ1Za6yrSNPp2Pw+mPO4IEHgRTnZVQmsN9F8BnT6yjlt2Pnr0vyubOGDPQl7/M8PensUS2
Uv4x1l3B3nGBC1tqCnU2dFkDkBXKTC6B7CtOUAfJB7mHTc/JaloaRD0+xzDLAp6vxcxphYPZHl4w
bM2DwjpMaXVk7kgIj+od6inys2AAQJiCh2Low8hPElvuQnBdB/tsOUXYpTPs93tiNlf5363ojav5
0c6ALB9Dof44ZU+H0VjdEZLy0wL94lTsjso/KpzcUFR7c+uoVFiT4tMWAuR5s5k9CY7fdE/E/9MQ
CKlCReDI6glAOynneAtrEzxEGuwv8OFWnLxhu+bg6B9ZyIahDT/g/1xGwSEWVNub4v4UlIFxtBSf
/cNLlq5oT5yso08Vn19SXZpIMK/E8+whaOeeHVwvBHSvt9E0+erd/k5hwFQxf4k/zzecVg7cIxFw
JStDFx3GTszh+kM2paf6z1L83Ga0LAcohPJsPDiwGIFCdZBsP1AgVcC+E5zKcrj3wxnsmfYwVQZe
DLAF+JmzrOuNtSxdODFBLLm0aYxzoGyaXs46D9EZMVM072InmbPp/J43rRHEsw/woFdXJovS69ri
UK0i8QBZr2/R6Nv4mPUZp7X6xFqF0ja67AeseR2+ufpEfi1enK6y7C3BBhW9QzrNPNS+rfn9dOrm
A1WDGCpwkB4p/va/fEji1dwsZR3LX4eQIC7lKzA0D+zquECsDwYJcqUrdjfNlKQIG/xJRitp0iGI
qtLrDPEyMTGSYZz3Pb72TssP7va1Zl45i+UVauYvxgBg1rIL0IHeLF6cgNpUKedUmw7wlPvZV3XC
n47/0762cqDjjL5ndUGQSPnZokm7uq14V0CqpfVrFVdistgSlpwohCqh2DX4cIviPEUYYjsPkR37
NDVU5WeQuqm/L1N8lW8Sb4DIlM4ttR5MY5XU5VcozZkDMpJ78VNAGbTTG2Z8O6vjTBq4oflo1hOA
uBZ8QBHe9M+z5KgdCRMj91uaLdfba2KmDgmIueVZ64ejA2p02fhH4dx+mpGLpCQ824MvXKNJOSUR
o8ATRzVdRId7njgNE+79y5syp9ZNMH3y/IzrFypaR2IbmKbw0+78QTsNpbm2Zgs2XDregv91qcBJ
Ud3LkVeFeH7TpC3kljrlhxdw3FPR94DnYDX8+ZjC9uxo8b+c2zpqatL7IM40V6m9fP9hBBLJ9lIy
5/P9KHIdbbI4n2T9JLY8VSwnGyT+CeOlQnHrSr4mZx8g2edi+OWqXk7WpjxsJNRfDOxa4QLhcElM
nM/WNE3HOU4+/jLc7LSZUAwYg4pZmUFdWCbkCD5DZH337C+kdJZHo5nZ0Xeq9MliiCNkK6N69vu+
xkiPw4ily9Wsb3vrwlJ7KtiEINm9yvHlsFVMmd6cy4Ctt5Rr27v2Em7ln7vIkBAw1YyfX6rRtVPw
9b1pXB7ozAM4b/rwFilWQtxeFQrIYDoc43BpTSmRgdA6nB3PMUQi48ntYr+Y7Fte144/09vWfx8V
96oK8wp/gFUWj4jgPvR128SC2XaD/zxUWQAEtHyX2UGVYJiusOkxTqWtW371+cj2M4p6Ro641z/3
sqtFmJJHWOjkFi68enas3cXCxoVnNkbEjzQzBD1+j86VcfB1BszMoKH0eh34aCS3SucmpciUXV7n
3f7L49+lK00fKHwD6e5JBDT70PcV79jvQ7c04S3LcXH5I+6qGm/5SIKX0/sdsrthIdTN15d/2hMD
TMBcjaBED6f1Wrpq6mTM815tOnoLQfWJFt3HZvvPbsCqCgKeBsv8q2gZNzRbKoTlDOyiO+HQCXJ2
Es2HZOUaOOFM+5Es9ULJHNLBdrquRDGtn9p1rybx72DokusanZZpSWT955lJIUh1Xpt2tf2hUGXu
qIxfCUM1quhQilWUue+afPJU7EsRwogVuZfTmA+E957z0Ksrf5rXadQKlorL19S4IUbYOEwMLrZ4
0TCqD2sDGv+j0JSwo8wvwsLhUS2KKM4nGTu869G9pTpa1FqMpHi1vj1sPCcfIEWE20A4zqDc1eq2
rVIeOhl/qppiOTnEVdSCdDAZA9eULH8FHYFVlXxCkCsTI1CGJjVc8VRq++c91YnMsMEyABBtj+BG
x6+nMynNo3l4fMdbZPxRPoj944LrKzfM+Ld20dA5NNDIIUb5OZufs8h4+jJO/c78a4RkjJcovZmo
GkQ5fl8rtISHd4+AKXZ/+62c4rMElwzNEAdFNhwXzawgxtZoBG23+8MlwF97eBMCYLROCgkKS4vW
BRw2XJAr2LBsTmN7uDb2dJ52cHMqVgBwZA5mZ0pUrLOw75WXUsV5wpgg7If7LRynsN2KivOEplqU
H/k4ZJknof9Sux/jKRHAjk9fQcZWmAiJkIfictXqAHOYx0/NxMtbXTbX5DpuvOOt2vE6qQO2WVrv
PYWbOBWZGAeQqf+mxDF3bUriFDpupcjMtFky8P2aZcU4XbdOKmL1q0KiAZbmecTwZ32kruNkOMUZ
6JcmrNhWLecw6yeSWYm8ildP4Yf8vGiA8Xmzj2ocfDLLT/zMTIFrst6AH/mKtt6EA3C4JsIpgvzk
urS6SAnwwK6WSqHT/Yoj1ro7fBE5iSeufXjKvJ14cHPMl4bMOIha/eKIgwJRc0u9OQVpBpVE0qP/
NUT51a8eUJ5R/sxJfmkOQz2UG1DMPbB7DEfmccz/pma21IY96PFkcE3XEvxPFc/ea8qJ/zXrg8o2
jekDxx1VvtI5JFoP6/QUGYIKzTYnt8wJD0VOxoG5U8uwE6Zh0TSLM016BoeFqpgvHJu7JhJ1FI8B
3CozbUdUnTP8aj7hE7G0oBWSFadVLfuoMwOxz0lSmud/WXkHEulwL0UD0WwNZDn2xtVU/Y7t6j1V
2p87jGUzownZdc9gXr1uB/IDrX/QdAsH1FWv7rSkJ2Dfjs7N+rd70fry862aq3y3umY867xV8IpC
8bmXH7YozcctGFen4K4kb33pHecYY8qwnYk4Dn/M1nhn5etD/cyc4zJtUgyxol4rPS17rQKX+ZMC
3weHVm+UsSIyRf8fdczIZZY1Uzy3z8acPo4Kz/sli2LPRpG3ZM/1XH870HAKe5/rzOqDng3ewgmU
V6e0Yc8hsB6G1y0YKjXNSvxCZ8ZICKtSIYf9VMdwgHPnMnU1GiC2oQBIL0/96g5MBV01iUzJNRrd
muRe5sNkfmDjPsdKwRvEPVTIEw01D3R/cHhtv1WHE4YBHQamH1R+7v5GiPt3JdGGJR0rYvwdfVdQ
bsq5NNbAzT5ALqUSuzyP92qJib5n4wV44GDfZJHEuhUQbo8Zb9gnZrxwEBwDRWYz8JU4AnB/xJDq
T6J+zeOvkQzGRhyzbSdCB75EgSDD7u4MyrBXRPtpCP8lrXYXCFvB8dTwUk9fYUWLBP4gtPPPgxOx
/8uPCZBG+UwyxgsCqi67WzTq/Q5GiwDum3Uynt1w30iOEymM59dIeq6wu7YbGuekVQsjElL0OHYN
BysGsz6Bzor7dHfZ0asvBxgOn2lC/oShbzDX7ULaBwTLADeinwyUB+8KcUxJzih8QxPqYbMJ26id
NK87HdINuD8PASbipV1aDSdsfolcdgNXnjAWeT0QpYRhlxM8zJThdutf5q8wg2UDYWAto2/huwG3
EnsQEF21jwuC+t9vGQ8xbJYyiDFjo+pq9AZHh2VysTcYnn1XjKQgUuu46SIyJTekkEN8lvK8HxuU
phwl5BKW5oPNd3LtlhEU7vdAiQEiNqR0Xyd1xzuzkU0apqXLMuDr90PeYwJ3Cf6pc7NBzGIWXO9f
9STkXrXi0wzs5lCD/zw8/jDfUwD5PaD5j/v1XOlKewjGyWZGzzjja3jhvfhzkZ6VlTdsKc6k4V8Q
1jXOpyFcoVen+L9heY1EyaVu0Is7BQehMY6GsOKJ09KKqS5jbNGrlcAETdIM+AomBv4qg2BhDD2n
kknSWPUm4Y7vFO2kocGecpBU8pn8SfWFee2R/kMO9UY4XRnNlD53Rrb1r7FsqT1EwEnAlV5Pkt6x
z9tYcO08TYADV2y/XHsHegGVPwa4vbVKKFX37/YxuJPKRCU6CwL9SR1x/Iblk/epZ9Oi92WWdXfe
lPVccDoch2ZBdHKdQILbPISnE8FAq8FbaVmMMlVQ0f6eRGhaJ/Rh/cFbFCelMMX9aouchEM3scRb
obY036FXiQuAeOTMv7g5/98ARHiGRJ50kIDT2Ui4MTHtMvzQwuTn0FSz+nOe8vV76e6JFG3fwcML
qn/kIPN3Frl4eo+AQqW0ArZ5xT9MY9vLYVn6+ohVMudz+d3YpZ5bjuegTk26wIeoUJIKyDRNzW/h
EB2CbFIMx39r7y7Bg11swdmHouaxqHYYqpx/traCXAVyRD+kAoriKAAPZ9kPpypqfFTadsgmNCKV
NZ/OrL0kXN2LNfXlQqXiaRKNvmASfvyukiMj6VRF17bXk3Poz9Hv2hQD9UsT+QWULu/0rOPcAErh
eoX+a+ffcFhajgjq+GeLrA+iKHUd061BVv9G6hb9W7t/nVPWFFi75rqI2avmjq/rk/dXRORYTKq0
VfdtylA8eMUCozA2P2MSE8Hn+XisvaU2eG6bp3WrHhoiCz304DogFV8GGr+O+xtIu3OYCHNQQwJw
hhUMAcHMFHr3TLsIIuRk2E/NbdhsuNkktq3RtYnXo7P3ftWpg4VG3ghm8cDg8miooRlGqeLJiZEC
F/yLJJe59kzrK8yk65qiUrhDMEVizZ1+D6DPNUyl9Gqd2Fq8x0dD6G4UkvzlVrOusLY2PtHCqCLC
FtLhMhHmD6c6ESbnGVj382JLhhl8bTXmtx7NBLMmf8nt3q8K36FXw6TNT1+8nGIee5Y3BCTZCzj5
3G8v33tBIK7ayKVs/m64Dq1nUmPnB8G3ORfrwU+d+n5wLb1Z4fSaLLglFZmMwTCQkYxyjpXLR3+V
EYib6+KxJt4Q9GUD5KOia2T+Acxc+TY30mbqFMvwswfDZEmMDu3gc39lHTPCnpjIMMEBwH5ffChc
nw782RpN2PNmN+wHNat1RhOgVsvtV3PmjJoR3VPgNgsZfZscnMbuDScbeUTc2EhhDGVOjFQZ2k7n
XTVVehppEa1kvn1f6GfQMRCGU6eT3UDRMlbaZTqruNGM+s4fjrnGGoQx7IzysPX4GY0K7fMbCZCp
cUtajYT2EaC80QBD63/8zvKO7sSjau+WVFiMxSunpGf0O9izhTF5h15Sz3OHsMbhaMx732g22TYk
YoQ+Fhfh1qVs6zODZfpgfv8axjf+6GL9/pfeQU61k3n5Ey+ZLy2BU9LgvQ6I87HqQN+paDxNJEFj
wL8kSmVuWPU8zHg6chJ6zOeXq36+149UkHDG0kB0PYYFje4t52EgxQRTtvbc+G3TPb5nA8XjfBc8
Z+KdwqHEcfIhWYw9cqU0Whds1X30XBaJ89WbpY+TQKLcDnyZqH3WEmUuJ2F/33fFMsuzLW1hUh4P
Ss+yIKoBsu83j8QvvewSSBKbC98+CYxt9R/FNn2ZLgBpaQpt07uESWFEC9sOUYi10tg+fOeFvQEE
cmsUKy8QYdBzx0SvcJL4N90THvY1yld3E6bgXWDRdVdaOwb+U51gcvzuRryQjiyH27txMrRh2vmO
iXV2pT1CzcnNPaGnlCNt7oCW1Y+1tTM4TL9bwROQy6o5BlY2UcHXYsBCyvNwIPtzcyICa0nDZLPz
T55VyJ1/xFHLXWGsQOsqrbVic6CT0OLMEnsYEW8y7zc/gihg25p5k8djIL3V9u4Njo1MFtG5Ygyz
HmumQD4R8zh28m0PTm2dYXbtGMhfPFfy2bQpDmC9mIAhf5UnTpbu2SP1/F0tN+qBGhgQRg1ODuXy
Ihkhl9ETlsmIjpyx45DACrz+6OorsrmGEZu6+BeLaf48fbU9GhbP0RAgEldLc+5bYuexOVn/YMCJ
KJv34qeGKVD/Zd2NAEPnotGKFc6aBJ8KU7yXqJKle3iLoBeoVnsadBuauDBeXFaSRQ9awVANzI/8
IiyOm5++2OFGXgrRwO0ojohzp2QwofVcHBxRrBeElEy/zvFGiNDLhI/rxZVRlJ/bFCRQpzZ8AjGd
gMgKxzkkLumbL7fnS8siEAT3lNbu40cjoq+ZEhiOeqOE1ghUoJDYA0cjtnRxuiraHGgCRe6HvwD/
UUdOr2qp4Fth0vtYQ6KtbfJcAMwAamYfHzkESW56l+SFJeWTu0JtuM13RZY104cM2Hc3oeOgHa53
DfuhOkNeyFWUyjOgF3VXZgTle/SabELtHpmEtJ/Z6VPyE4xVjBAL7dY0O5TYatRJx8pIM29froUp
i8T0mf1cNSe/zOfb0JIp9P8rkgUGmIxEX47SjsHZfYBdxXR83mA1Q78IJGzSWUM1Q94ApUQaukQY
Rn1+3PdLAbY6vNjVQkSMpxCrF5QCGk68FwII7hhRTJ9UKWpaerttq7fMsY5we7CzYm1MK4d1xS5L
ZJb+JnvDik9RfDfV6/VRKmgbWq6Y2kPblly5cWtYjr3PnEkZ706c3SBfXikeAyavkcZom3Tq/V0T
NV/SxNkoWDOHK8qBVyWoKRdtvJ503nbQN/Lw6tHomR4U7JoM9Et28mD1xmeq7Wd66l1IQaJ7Bd7d
7612i7K3tF1DPr5Fy+jmfLXuIa8oRdAsDmwMKEb0w9SrzTMu4DxhwZ4xUaC4wHS/K7O1Gkjb1nhw
87eaUgXweAQg+TngTl0ahAT5JYmQxLs4jp7dzzyN1JLym86SIXcdE969r2GugDTwLTIR+f6jD5Hi
/GZdinyvN7t10cuYsKMRrq2nXgfBjYe3Xk3Dc5kuCnsmYI68Lf1VGaZbblbd7gvKmJqzRERMlCkn
ilaSVN3K7hWvRCjO3t7GYzMQiuqSUyxwUFFgil/3mmmP2fUbkOQp6NhKTERU3mHkebsapDqedYzU
yhDF0vn92wxHCiEe+8jBhw8mAQ66xEywsivk06UTgikF2iFZUaDACsdhTBz3xQn6Iv9PPZAUSfUT
ERdpUxtUuaK5Ev20KP82ir1LVpLtzIBpPUpCYzC65jP7LzhRyZfzR70ZaUuZJQN9qK/t2Vtq9hSJ
amHNE2qZ/f02nNad6TIRmevyXJE0Rba/AHTc2BhN9tGlN+K0k60I1rF7DpKL47oaobN6bv5BDUMn
1PW21h9817na5dL9CVtBRy32mjfsV3vYufBokVyUiK16Orq6kxjfMAlkTIp1BALe+Vzdg/GSDOBp
I6nOTXlq/yADpVXoO4Fev3kZg1rAefVuaSBY5/DjeOSs0JLCHSA3+MRJ6GkeNyvubv9lEfV7e966
jYJ/RqX4QavSsnyE9+gf4NtjIWl7m+fNZJWmgGKLyqGyA5F/gIpvMXeBeQ/N3UThI+CHBbYXnr8K
66/NS8Zsu8SgvqRl4OdQIsgBJktKfDOygOItdrOWtWc6c+SayuJnX6lEWdHOoQFyelV+xPaY/2BW
w+A1i0YaFaCL997m29aCF8hPXzDtvZhkMnRCd9vVcPnsBo24v730lfpeASOAVivtl6XOFkvXCZWS
H7aGQlXITIvewShptog9fswjsPiri/m0gVTsbyzvuKzJEFUG3RDfag9tgUwIjLjK15JXZLTEG1Zc
/nUEvjWn0mvvO7znyMhnrrJxnLl+XcV2WbQs0oD2NdYtLKJi7Z597A5rp2OFjvsjehzQtF5W1lIX
l8YVhWDxno9wZCQvo/3I372OsXshHkVN0h8W1/5+1sRZLMuk5SPy3sxj1+9eIAB8nVc+6X74HoBm
yXrnoSYVnme7uLJsXQfQJlJbfMUcZ8iqeGXYJc6Pv6/QrhKz41oXEbP33iNJWoxiGvJoG0aZYQqi
Le4BQb6w5L8w3XRNC4Mkt/0i1Tn0uVhx5WHERRpFxGiDPlY4gm/A5YMw/uPl+BbcmtNiuy0XkMqf
AkhAnEE8jb47bKkr7nV+wMEpbNx7JD3jB6ukrPby1wdSVJBEvxnPYvtYXvfpJvgEmsRoR3hK1WfM
dAEjM9k9XOA6ER8HJB2RH6i7D2DACjrH+H13j5MwQuUHcbMeBe1qhNAZYDeEuBROJOUM7xWLtutz
Iyc0Ww3LkPS+t4VcYu/5BlGPuo+RVYtt4+T12dRAaz+uu9kVflHkKNnfHqrfplRde2kZe9Xcusm0
uiqqwePgethI+tKCZzGIDxmUx7QpUHKg5dA4kbYZhR3GOCQFoe71ccfTIpzsexdXA6uS/bn6hMyM
U8mvWs66LJkaiSHbhoOuQEZHkk/VMoNRli2r2d3RyeqxECTn0sxoCRiltQjhrxlacETE5ZFWM2MD
6FKuGWZwDeQzDVG64715/6N7SP6KyYoNTZeS2FmK7TEIEAR+e0FMpbd0NfG3Ni1UWZTzM322Z4v3
DRDEh65jnoH0fCqlGz9dA1yUqpWbytm0s852/jEfF5vimM66AepJ9XbNzn1O7O+MET+SBNNR4sQp
tS5BMLyyC4LVD3xk02i/xK5+I1x/la5bohdFFdViLvaNktCOXQgNgUSQRMUppQBMpxaWYt0XhMJJ
6OThwiIZrvPkxYTP+Hd8gmiMFJicWXdykDzZSNH3bgnfAPtWxuJwKceJSBtRL40d8pgUKpph0iqC
EEUuQ4Wgp+ezUbk/gq1wA9fJqPaLokd/3hT+VdqCklrewU3sz+owyAEWURTq4keU9QVRhcey7fE7
aosJEP2rdGlX9r0XOX20ISEhrUHi7xOOWMCI6KdurMQFiyWJM5CkcRcB+Vbaj/YQy5kA8gMG7709
z5gLh9iNfk9ATBvDZHJJbYTwlXR7QtVwdzndJWaqJPMR5xpigqrJq9lbZMfdT7tjLqNQFOXvUZe/
3ZXUzf6f2bt+Oi9IQYSN1v1pf3yWWSMl9OPgn4DNAI56imDlyBjkMDpf5ARepSKdmATZr2R0292w
k6zy3AIqDLygUs9n1yFKINE/bJDmdNjnAu7RgDSQ6jGE1Dp3As+xeK7H5FE3kpzbx7IdyVuVT0EW
EBOl1VAn2bLaHZdsmCq5uScIRVOiRjn5BECLeKaXYh2WfO9p8h1Kw2NZGHaqraMZmKfo4J1Xl4I3
b5Y8o0JCqd5QzufWUrUmDVOD0TUyGx3L1oPO0l2JC+tQxP4XooaZi0Ph/zXPFsR0qmQnLfG/g5nI
nBcKAlcu0sOO1GjZyAbq+LSTlwmO026SZaAjp/VNusfq6JoktSrFQJbmfxAyVkVfuLUpC5h9jAfT
R8vpgwopnvRaYC8HPqLYDhPvWULCUn4yJR4/WT9hgpXWqIyo15XaWsi1CfmTNCa5yt+haiRqqqTd
KeL/LeVg2AyrEYankjyG8sivVHzlngDUs5X4PyX2QZBb3xRG7jVAhm1pBC2lSGjrHAZcHamhcJOU
WMix1igAZpENVJm3HUJZQ6xNk2NggdGMnwKcfkjnVE1Suhve9NA7hMaCKSfsLgZCv4B6VTfxnxam
zkFGih8IcyTu1ODDUzzGcQKp7/IFKKghY8RaecUsICDOg5UXyddB4lW48yoVyRQOVV+t3JDGkfGf
RrOV3o3/wWnRHjO2ODye8f0qbSR3ksvfNC6seDtlzInDd5mgrUDyRGl7Q4Y2YtoR4fhyv6rE8Mg0
taTVM0FezDXicumWFYm8hQEjupH8Qs6IqBJ/FcJOzuP7+huh1wEb62UzZJjdI8MUhNlQ2+EJjLVw
DYFWf1tVdQEeUdm7K3NKs7zVaZzxhEAkkrhPgSclqorK219pXcs/0ZRWT/901sPOatCXxlnMEuWy
6BGGjTSrp8Nky3em8r8pOxpWCSJtZ5Rl6DWZGcsfs8YJ4ttbvPzneanu+5xB4QiOh6pw77kBvcUp
AvvFLP48AGyIbZOg+DaeO8NsiYeT2J/4hM8BeE6at/Xx4dDFzMWuQ8S7oIM5y5fwAp4dwYuwSXC7
ZB+AiLgMbsz2LpJfTWftUuXiw28ZKth56EnkfwVjth02Ggd56lCJ4pjYUxlFVqZIp1viMijcd319
3D2ChpeMqVA6rVyhmG0SKkQonTWXY9JpJlJ6yXnQxcAAm0NCCAodZlX+KuQWFld6afYRSeTZTbfr
bAViGVFOTdiXXwywtoIvlNxqetkph0+gBsnS809c6XlywYgKH0JA8gWwDAmX0ug2bwazEJwxdlJr
mteNnAqR2/8FsyqFRUQBCdBujq0pjZ8T0ynvQGkwELsF8cY9/G4/JaytC0ARpwHXRrngDrxN7aaw
u9YVXL+iiOYbClTEt3HJcUZivhgw/RS06e0cbGDZKJ91hGkXLCfx/UUOLQr4K2BZXgQdz6gfFj+A
FsWkIC0p4zG3zP78YBGiHy+WWag1bIkpbumGCCTS+ajzF6i2JRMouEtTXE79ITrXNECVKHdMib4T
BqlTHsM8fYvtsY+uN8gcDRUjk5kkcuTUbzVI6Ya2oirRWouji2F/CuGslmS2TiXQidH6H28xpELw
8h3b4tYyk2lGzwSTI7g8K35kzhhJb0GIbvS5GFTT8SfRpmpmArkx3GQ7aeDwDuDyKsYe8GzicH6M
76to9kSs9q5k0yHzz+aVvVYBOdwsw3ZSSCihwU9d+7x9YnHrysQg+VH+jgBVPuw2G1zhGW9RJfOK
pwAaFQWNqqENu6v5oc5qlEA3z7Y0syxtRFiZmFCf19DKIUpTvu8aukO4j7RwT5D2RR3e5m/ipucY
okGkyxyHt6BVrhyrqBXk+hGYRtrr6rObe2xzkx8BvP0Yej53REboZLk0py4jQRMSyCUESb1U1cFI
fI0+8O06ON9Ia8FQsGfQXkVb9JZcNJaHcBuOISuIC9lG9QiBG4UcTY3mAw2DdFAzGj4G5QjXKkrE
yLu8q5gQdiIVb35iHEdcmMhlaPytAh4/pB+AqjQUhm1YZLhOw9IkWbG89WBNnIAK9IIG3UMHvNZt
GLOBpeYdcBspbkvwTR0Sn/6oSEYTfKHnlS+a9lWNkZHVBxFs2WTyapiiqdD+jiO5A40CuJK9OD+9
luMjnD1HMLbM0RqY/gpca5S7AB6TsIKlHZ+bCW68KFCgchtY6S0U6pMKVhtnGwCHIedF2F3zuFd8
8a5D+Gvvk4OuZ5tLevS4ZSGykznf6yb6SaZp7agKiNpr0W8WXk26tQIMRk2O4ytquqcYsJcy4N72
iBnm4cLVSPxQOihMDvXlZd0T6gWsucKVa9cLKRS6xMw0a7Vbky0Dzzlb0DyjwObxOOu6t2pViNOI
aq4Z8bp1/zpdHuvVGCoQyj7ZUo+AUoM6yNGIIi/3zF7W6fVcv9THLS6x6w002SCTnCLduIYJUctl
vMkHXNYCwOYWMmvDIGo/DeVT5Hs/djS9B2qrws7Bv5/nqwn3ySNaJP0CgORB8gIoN4o/OCkUyyLd
pLAY2PTHmXp8CmBdaizM5B1P9wtWropvPtb81WXxcxK9yfHE2XYT1nkXawxqbI7R3/ebaoN1Ss1g
Z6gIT+DSsOAsCrtRTMa9R0+q7Vjg94OVDLJhvOhzxdP3SEVbf/HWDdjCrKj2VpXsCqvIoriJjBfU
ln74BfLpMjcQDunKGnRU7quKmrRqAxR9Ya087zWekqWWhDwaNg0XJIhZWNRzvUd4W3DiH8BQpseL
x5WMAEsQKLaU7cUm8FglHl3zavtVuoZzdwbvVJ+rxSvf29YXGT//rz0aMGdswm517oXDrXoZnAFm
PMkFI0PcUite6ZE7mufFz6m1p0lGAWKuWRDWVDi1pOKlf89FOF+A/4fG/Ud/f9FEG/XXBxq0pC+M
Wwl3WSF8FHtB2+/TQmejmB1pSuiKiWPP+68EtRXiWlPgExqhfWSfavhS50zoeceYjS31x09eYMIK
2w3NVRsVWup6TUdgXGL0HUWOqWrK+72tduLkm27M+S7YVqMMTgFfpankY1cqAEED/SmrGnHq69Oz
glBmH3htCHcCaDRU8cxLidyfWPyiZpFAClQqQkNHf1UJFG1mK2UBoAPTwpBMNFWPzu21YUCAqiC1
5AiM2rUMRh574rTf59f5sjYBA1dmxv8ZOr4VAr1Pbe9JpvptxF9pXexFjgnF6aYdwvOAIRajWk2K
Le1Ea4GnNhlr+VWWEKow1XWflSJtOzI7+7iDhM2K2mQ6l1VsKwCB50ZnkBneTRx/eLQlTJxp5eq2
4dw7wT0TQ3sSrsHMLg8xQTFYhTByDGdDL/nCECKRTlOg7+cvGfgonqKt/SddlP4zWCCl0zcfZ0OX
NSiL1P/kB2T/ozM3oMtGKeO9PK2Jxw8khPZ68aUrIPveK/HYZ4l20lLqoG8g/dj+Ev5ISWlKk7gw
7oDPvwWJ+yY6n2cJnKxmdQEr0rhpEi1Jv3rC4UBYhqmkBr9A8j+iJZXXqj/Em0QoFqZZdHezytCm
ECsSgTl+42IMIuVIP4T+k4DcdoRYzFJGUdGwu0/IxVRNpb2qk8HfskCpp7/zMzaolALkfR8Mlj0F
ShtWL4Laa2w9RUivMcSU05yG6VnuBWWRdc6bmEmSw+249btuga3Iq3pwl3+rXltH4/e7i3KT8tXa
Stnc7MzpNpEohLojmgczRQJYGrRkm1ehcwZ+2Ooa2NedjRNk/8TiDcUHKwcIBo7x5zS25fZBbScP
VViwBLffb1N8Bgisn5+d9taLWJ0k9D4rm9AWlgVrHxYEfwhbi+sh0TOjmwlQLWRKEdRNzc8C0wde
hp8bsMq4Mlqsaxtw0OU0koUEtFvJGAA5uwx08SRYeDwmoMGFty0EtxIgefyT2OP6LLlSsClvR+m/
P3gWq/PP6H9NVj0RGWNPFzxsW4+dEfUbU01f+Godts/WuCyHuYumj6t7SkJZXQYQ/0tNIDbL7jJP
/xkdhKMi+LW5W5THmNIFBzddXtYW/k3dh3SaJf6RLyWck+2zXzxSQhvO1G8+H0Iio4xfm+D/2Gss
RuiHsWAsvUGM3qUpWtmzKwUTjCZVyukAvOs8iDxeRS0AcfL5wS2xl0X3GY+2rVrA5nIz7IX7KEZ9
4+K9chi7DK+ynZn42AYUunAnXjVxFYKtb8yyikvjBF8fcdy84Nv4Dtu126g0Bb4mq3WvWRkRInu1
h5Bn84lNkjvbhl3sCUIir5L9q+WMNHQxRcBv5Z+zYgVskgAL2l96USc0tgXadATTurQYMh061bnf
ePzIdQqjeruNuf5HuMhVrGeRN88k3WS4MOSYZkkwh3B/6bkNAQncMst/N4+g+AWXP8Po7hmxcn7O
rvZ8EfDU6xjq5W2+GtobTKOBIWzWlw/L9rBUmb285uWbUx81WAdh07dGt3S/cIWVaYj8w8Gg98MU
/KzUgX6eX02+Nu9zzyj0ChluDY0y79dtL/BrWCjv3rFxesAJDnbEWaZUkOWtD3vWI0gCStaySVEG
Bte9fpHikrkEjA/DsqmUu1Qk1fkES1LCej1o1dwJrSZqy878xQrZE75u/uaxumN+4KyvKZv02pfO
vy4mCCiqkLF41D9ovc6qEf8b/IEWkASIexmt5xISz+XaxPvpFJsMYlfqHIsbra16KBZ6L5D48Vh2
TPQCiyGl879482f68EjyMmO0KAnFUgCKQGJzx6ExQBMKZHkj848t5oF/XIWbNEu3+53iLrCrjgLw
gS2I5/6NGe8+huazjbDly7let0J4NAxMk6nmhiyRZ6xuOStjHz+BWDIrlnpKaEssV9tBkjyVT5RT
FyvCmMSgCzJltgLgK7D+mGql0fed+CAb1LOzQPryRBIyTnHLcV8ZpWWSmFtIDoblGCDSGrI+TBEr
Lh4U4Jrvrho4hBDU6CrlCN9wCfLmjkZDxoOuAuYzmgq3qw9tByEfdDRiGeCq5A9Qdjo0yiz4kfsJ
9AfRphkmqQ9pC+gdbwJkZnz5O0FCq6uTKTxP4MyrazHqswOuNEht0q1B57XEdvnwrTSlS5Hs+Q3z
W7LLZWItZpLErd31UOHSRNjzOj9SMsTjjwWt3i+t7SCKyOQ7GSlQ9H9BJ+J9BUAzQOqgFcgd6zbq
y/xIctKtNu+1P/+IgojnsBLfj0/sKSQNlwY6SfgvXM3ADS6M9/V6genOsNZZbKyHNQb9rbXSh1eb
aGxtUhWQn7itJRb6i0v2jduVwP/ODo+QVuBscRmpE3TpXE1FtczAKdJUNjcU/l/MqP0LWoF6ep42
AAbVs5cmp8ivzSgbHSPhjVLUACDdz36opUjwk48IBtyxFfrmlwu3cu7RLGAljPBuh1cEJ6LJy3YS
bpt+jtjy3SoS2/aGBKcXqrnoR0bH9qX0AYjiZzAhckM7gZCtjWsja8XppIzk90fheS2RbbaWdn15
xNBSwWSJTnYf96q9IO9yVyfrVfA1nXDNJWNpm2A/n+QsxH3gRszw1Xpp40OH+QblN32lexp9soCR
qpp7wb8ThuS4JuMZ6yjTJfVIL1OtH29Cf3BifgFomnQ1vawyAjqPGzC4TX2LLzdaLnZ5EpCQZnpc
mYzxcPVaUyCLj2e1fYSqCdTuF+bdr+9SYY+RXD/pwHG2kQraUzozmZ26eAsOJJN7fRaFg6NiXeub
9o8baRF/CZLu3uOW8Df/F+G4ojyyVNfxYS78sKfA6sdfldBuNH4srRg9tVCYsG1LtHlycngWCslU
UTT8m9Ru+Cm2Z/SQM7/dL5q8OpmJbU2HwesRjiHTzb78UvpDBbvCy11cbPVzEoIaNa/CWQFf6lZs
AhC/Uwx6QKo+B8k7OoUkxgc69jw1nSvrfjGnHCn1eV/1LgjWRvXbE/P2nlxPuQ5wWkEOykfMrxcX
nythnLqPHQOmkOZ1peXvCpwBh19JGFZuFqlf8+QKoM725sSqmM7bOje6/Zy+dU4JaKRTg0Xjl+xP
TQvgyb8XlR9/BddJXnKRk7KBMij7Gg7qSgVAeRjpkEVgyIQuxrj4vRWcfPghmbJNVPmMIwkh+cPY
vWf0fLpj7DfpImodVe3ewFN6j/i/u/1eLDejVABqrh3cxvmmwBJsF1/w/VaJSC5Vk64FMrni0PVv
xQDpgMDPAaxkIhJ6izbeuKv5EKZTSupBp2ng2seDHZYQJCO+LsJXilx1OmAsYC2BjcGYprCy6c2Z
VGKCU+MLv0sPaK6+jceiBeaWoRhyx++P8fp8qBhvYGgMICCrPtNFMQjT2buAoB2dpO5CMiuE0N6F
5TMXqPjgpHbq7+M3odE4od4HIsmCSM5l3cUGYK9UtXtDK0ui896aahw56EhDfrvrGav8nVrHmWN0
jYqtLdW3P5Qd1zIGdecSltddCeHlD2JXqSO4qwpa/PmNnC7pMLC/XH4wWLqSoCO7gxolg4ziIj0E
4a2/oSdLfR0HVosDwOnhk/pMhz3lcW4lBTD1YMbOY2nh25p5uE2vBhqZwlxQ4DSOa74+EcRGtZN4
nGS4AwRcAae1q9bphjQfM+BhliKCoH1DCFlRWCvMSOYynMPQer5jfTk5/kzElbOuswUhnhiQkT2l
L+xwZlNvLIwmyIYtn06frnOHNUFzKGYlQ1A0bK9go8eL3JkBvcFnoLIHKjKtzdeSA4JINQoB58eD
hiPVn6uoQYDCbeDnpS9+8NjxYG/2D3hJtNou1tCieNZz3gRUMaZcaJav8Z2rDx1j2ehfTXYSfxsv
eIQPFRj6uQoTAN3e5oCsRsR6xeYyNrYz7W2gqbOQjrlpFWYi1nNoI0g9QUMMHEOXkcee/kcdQh5Q
b22G+sHzLEE8V+CsdMuEmenBCcwTpyGLTaUlruarqdmXYEdUhB5wEk7iG6YLsVxQXcJH3qWIOSJW
vwltnARb9eeqg1w+ZDmgd7eNtOj1JGESg+tm9K/8RzJ5mU2uWN/42SYAtdbyGPb9hIPozft0CEnj
wYnr5RGeTKjgZneaXuUBpV7iCddAa8xzlxV8TwJjTbXmx/SL9hdt67hsKn4lHGsSlCoOGDvC/0TV
4P1ZZjqDnCv9pq34X7pjtOKrxh2UNNq+bik+TBViMuw3nliOEW7MqM/qu8+PJRiH9kvNz33mXt/L
ATN1NNq+lWS7Ki+wG+vzDwXBKhPQVb9hBfTh0E4815nEzqBy5PMNt32UElNhJz1beeRnisUKgYUZ
Emag5GmjZL+XN+DFE/YvEpAtrBfkY9bR6KbVhfNEs0scgAVOn4cUzr6sRZzXVnCq2T2XegJ+3AE8
gmWyRwAfDwHg9uTdiNTxhYp/lKjHkaOKmPGbEiSUgiZY7K3/Kg5ecakG+Y4IxxvcuWjDa8zVm66C
uWARC0eKevJ0/uOnILx3Ywut9PG6mcAJYA0xHz/V9eCTguGJojx58C0aNaHLWhdaPWpHB8C28qRK
cZZtKzUyNUun3I2iKhb9IxARh5ZNxuNRo9+YhTrVT3cwRZhFFgRT+6wL6M8hvt7ASvKlcd5vrOAg
keOfK3AbAcR7aSahnC/7exyMzqOfznPh/rcXcdnmRbG7fDiZZfBlX2W5JvJvcl57skrqD+oNNw+E
95KiwIlh7dFxhvvlGadjameToc+qmOqoRyTkbGaDF9SJkvrim9MPWd4CdAcRFE7KqWESRbYtvjXn
7WZs6ySrLHp/c13fT3EdjkCZiKrDXLq9qrIWhjpwe+y/pdoxZKpfdHt4btED1yj1VvxE4mvpFZNx
iWTQc9BmeQnKZHn/mJM47vsxkQ9TO/jvx9Z4TU6Yq2yb/jw5HJ44rBT+lLG2vepY4EBruTKsed/T
QNwmn7nniV+8uNusj/I7dd8g5xtpe2SK6GTtXjrxr7k/Zv/OvThDdfVl6nAg51NINFjVOWJUSPOQ
SufAJwmclVDyYP44BxvrmasPe9SOdNMHyp7kb39fEH2lQXyezeOvO6hXbxSGAqXmZfwtsQzQ/XlE
dOfbl0JbmXmpPK0wEcK1QZADvIZLgG0ZCNF6bGtuixz5lS82ORiNKCD75jr5gUf/xOuI3aIUSDtv
4QD2owGB+ilRJhnEpTJT/iaO4YOX05EZK+6wTojStYsUhfYbI4j7rLETDo6aA9Sl4ykgN/rY566m
ABR6r5WuckXhu+zCiGfnb38wF13Ad1AmQMprbd46XcBaaZk1NZ/HB8/1tCGW0eBn0NKmS4IZu7ua
PkmJCF5XToUL2nC5NCabrUlNL9dXRX3QKQ3/c7HFKnsThRSuslsBkBRZBBfnsRI86T4uOFx9kbQA
7ai9Rk08LzeoKwJ2P062RBBgN0frENU7N8VztBWpWBlls8xAxQFU3fL48GxZLNeoEAk1vyb27UQE
/hn85FvnC7kUER0WXOpg0Kzwl6W8GrdnblGpe4BnqhCh9DMe6zbDXYtWLnjj/UZXXwNVIsG0uAm+
x5xNt9A00iL9eDrmuVjXYm9rGgVwO0SAnGu7VRi/cn32s3ROBnZyrlKQqvI+7/EnpGs9hrk6iqKO
+DIJLOZxLbQ5pHkYvvd/xZf0QUBEtrXPy13cdn1X3hoTaoYLegLbYxSisx8i3PbAUebYdZuJ9vxN
7B64V2bHQHSnjLigCyE8CeJ1XjdwKr4Vavjxu5tu+TA2qxmSu7K4X5tL30Oyzk7coWUTdUIU+H2g
qVeTLM6u/HTMZo3YOsF4vDPu+MjixT9D5FyIT3ognibzE3TLaoea5ggiyfGcgBsRbpEBNnaRgqjQ
8vrLxEzobfADNH/vqD+w4FFEcv1tFFi0uQOfb+/hWNheZfi4SdD29/aWaIYi1WI5Vw7xz7NefOwT
24AEYn3wdRe5G1NlE7bIATwxcoihAFMI6bOyzG4EwcTAA4GEPeVafsbszIuxqRycCMiN7HShCOOI
BNGOuqK5cQG9J0z09s4Yr8qG+4ui454yMrp9gRo1ACzhOdpA7b4SMnpQ8mGEagpN2SRyGJtKLMr/
Ki9TC1MMgilJpc0hNBulGOjwaTsW7VibKrat+qkN09LPMnYMviY1g5FgaOWRR2Xe1mzXyATIOkww
G9oV47iZ6IKbix+AkX2VvwKc6Vht1FJlS0rpK/Io9ooLyubteXUbAbEJOynf6Bn6fseDIoP6Wlwp
JgNN4MDJQ2FQieP0ezXso1LK4KStco+wfr1bLdi0nPt5B7PDyV/SHZECU5oKhugKrneP9W82n9fY
IRQ8z6YIG/TjQBKY6X7XCCLEJM35N9a/2vcBlcs1frxQmxG5pWr2Dl4Y7XPtsBkffOrzbZHvHXB8
AY3ozyhNCyYmApX4Ksmi3/R0JMlzwixGbDRuwwF20xE6g2JfxDi876CtFfh+pvk9yJkd9VkoR6fM
pRRtRP5zf/KRIZWSFUo8hrL4Pu32PQVioaBM3wKclVXNAcgiH0+/IjPxcpQdjPrt2+qrYdIGPQ2m
2dhczvowsfh79SO20wF9r7uBZGir3/9NxOrfvNHAhbxqRo/QW0ovE+9cwSfsPGFZyFMRixTJKL1q
82l9iJALvKlH1js5hYXu4qIM1VLN1YaP/yD4qm75MJO5YgsifxgHnTopRRsP5sMaVWTbEu6+PNp8
RAB4Uek2z7lLdBY4ptIdRrWUcgBmZI0ybZBgCUmqP3r2kZDBzxDSgyRNH8f8IBRHlLDe6p/Hf5se
WrpE4ral8+CdfXOZeSP/fdSaZ9F0nrEjoUBPCBKAPyV0maCMnupizu9GJiuUyb1/CguUlOdF/w7t
zk3S/MBDQzWBDbLvRjPNM97NkOxN8cRWnOuwjS02WaA0NeBxcAxA3l7Udrl+xS4UvIG1IElTq6x2
iUan3yr2TaDm3lyQKOGheokUzMEyJIuSjFBLamP6096FgCnT9eFN0BcTlc0hvZWWnPHjRez2e1kl
KvZWFXY0kYeKkWTmkjeDi9E+CCOeNbnpTssDf8krqHV4N688cwvxyJPYauTt7D9wPv6GkVgsGo3t
fWvG7aGzInBTW41v6QUHroCb5MN91THw0SphwxWxpS72phgCGzFK4RGbBmlJe8sCKj7iiLQWY9bk
2JwtDbKGMxofa1oCVKyjXxX5gTGSrjTdjRMYURE7fQysKwEWKTA7vk/rRAkxCo+jg/eOoOTsg11f
Qqi1c2r7uTFITr8kfzimqYQ17wPdEhJlOwq+qF12kYkV0grfzifRprDPLWtmDGz2pEVM6cdzr7S6
5Utuc7AH+IMiT7CmGokPe3By5QyruIawqH/bK5nOnKgKIxMyP+xQfcF/lON7ZYWFYE/DfkPo+Lq9
GvGsAI6/H5vlFoV4sCHikg2JaUtBMWQczjB2VwKepLgxBIPrI5GySe5aRhTuzbXZGFKXQN/FAgMn
jQdZxVdBqgOfGZBpKe6kbzd8OMKDNvmSjVyYQl7+LiERPaQpYo8VE1Vqdk46lrzdqDceLeCPKPqe
F429WKOc0H5JrLHL5TuYg5bt70wiUZRc7X/exiKpfaYVky2BXjXxzk81co7+Fzkf7HogC4mrqUSm
FuhdYACVPWKtMTIB90/Xo6PTNcg54J2WWmab3EFzQ0YpoZKGzjeWwAD7NVA3vpKLn/95wefoyY9C
ZqwIzwNpfU10E/EhG1uE59QGqzZT2/JTDhDN7NBtkxJu0wA8ot/qy38fkpD7tZb82tVvBDbkMGP0
4kf56BG1tlKW18nJR43ParRLMfSPfjwNQOXajbQgQkzTdW+a1Triax4J0z4a1BfxtR9QRKNVSeke
yQbzHomvPkQ8DM84Bwjl074AqHHwCLauCbLeU3hZPg/rc0tk2+hRXCb+wPVtj31UzLoUSgrwqcCL
7He5ljBJulPtbnoCrk2gW6kkZ/RL8/zjHAJY1VU9roIR4oE/kjybrZlxWRXWVXfTokZKve/+GWhU
P5Au3eoWPIRtT3MBO0FVPVAnmceX7dgGxNRwprizeL27lPXuA06PSk80OrqgnCg746j1Fi9choh1
zcqMJFJ9aM90bcR0jQURjNLymtqd4pAOlL0YHA+Iftsb2sWtR1pQw9tiqflqx5KgUsgwG8RS4ofd
vBu28rXOzuJhCuM+TzO6Q3B26jDreoneDnX+XjuVPqLW+yrvF8rehUEu/QPmtN/TurjOhUiOWqDN
CcmF9cSp4YL48n8rCLaXYs74c6Tk0uOD+wLYiSFAQeZgYHW0NhFOy3M9MXyz92xCpC90TgCfiKOd
LH/M2aA2PhflbG2HqqNDFgwabKx/8vlpaUvKPhdfe2Xni7tmonPyrPoix7W9Ry2M/6hqC/m5lctN
f4+2eIAqu2xnKdOg4ikDt5j6BdWWUXqFRsLnvmLdzZOhVA4lHSM/a358VM1luf/NjD7NiVw6MOc2
JJo1KBOWEPYPCGg0q174iHfuMIBxmaTsDhPRQZhwmgCBhQGkSo5nl4lXuzCP6kQIOCT+c5B7cyq9
1ItwTT1ooxwFPEmA6GTWreCIficzpMdWVmiABC9ObOedmi3o/9JnR1UWimjtPliuQY/NE02Oq/B5
7tVLMRm8WvPXQt97QRIEGQrexjOq/0vq86ZWfVFOC/Ueuis1ex1pmMH3hRIxu1gyjO24dI7/oJAN
+5FX7eCCj0Efv28autEYQRQc0ThDNtx0iYJUXJL54VkP9c6J9Bj44ffJ9TSrwNOS4KLsNmgbdQ6h
Dl21eCzWZ4qOrFOCKWB1QaHzMIthe6vZIHRx/3hdVyLOUHXvVg9ttn2FK3rKeVvxZPkEaWpywLxf
0/HEhs0SwphOUeMY1zWWrShZfD+FnWWIV3xu41HrMT8DdvEkdXBMA140TGW3mC71RzBsvSq41RZc
qRwj5y2zFiGhNIxDEcDDjvqYJgiJZrXHhhdwhPOZUyPo1vfCeRznYZZfcXg/DptL7/jy5OMeIUZB
IriOCu/6IQ1m2kL3zsb0dPvBDAkUS5DADFPwO6f714C3Z7BLQMwBtTN7tGQTdgscaZc9pTG/nLJM
Rn1gXrGniq6j0HpVHbK9XBnljJS6J/cTY66yER5LNvFzn6SeK4Noah+sJgxRrv4/xddgGVXXShs5
tYCH44OA07TaUVjJSdxhIinGcysLolVhf/PtRGKdKCOCLhg6aNiYd/QBzzubrgwfG47/QdKzGFue
3hq0pln0/7vphx+YUIRJjl8jp5ieeMa2FBB9k6GY0zT4lwkhTzvvQz5Rlp/Vz+BaJZz2U1Wo0d3a
JB082qv4r995JkcedkWIMyH/4Ic2cE9N3YZty/FcWNvmjfKMEdnn1Pf+gRuYJvttNDZxI8pKaPbC
ycjkxLjgIsqeV4etdGCBZHCW3QlwV93M75cMeCnHZz8ej86Wa+t3g0Rq3F1zanYIKTNYXRtB1K4C
AedBs2IryOFml7yz1dvh6BGWB+XUp1vlPMYJ9yyzcPAsD8xXB0FEL3oyXWMtv2BtUxRoqDnLcUvA
6PRIW0RK+kkLV852wDCOiZCuBJY/HOvEB3KRJSZl5CTNsKne/wWMdY63EwJF0NJ+4TOc1tEiovnz
I9cMC4yUUu1u12hsKVNFlHkrB0Fycawt88bAQBfxUO0kVzkfSPLO/fHPS1xFehjeXuyKtW6MNpTa
+3c6MbFGZUyFX9MV//2FXTRs2Ax0D8a9U1hifSszHB6YVUps5XNPLaDLSt9bFtUyC9t5UevduEj+
LtMkNj07xdoz7kDEHCFlKuVBpgPyXjb7S79V5MJnui7YpeHMzqGzo9aBRlGLd0LolsZJLBae1dnr
OK34B3Rwer8zB4weRgT32SD+4lJ0EWgKlsbcvrxLM7LdI/HwMFBHbuHTy/YecThoCDHtHMbeenFq
d3GhYbWYnYVB673NflRdMJY8blt8h1bcIQPZwaNTCxja8DCsSEucz1koD/J4uDWV8+YratetyYkR
Bdc+izcMYWCuk4/XKuzVbFQsNbnMR68pCwxjM4lT3GRvrMl/JC6XJnes7hoTtW0mD0JR8IIvf6Yd
Qh4CneJ9xoUBuNuND3DCOy9RN0qjozd8fEoFXQJya6VRAWByMN53g7N+4ZLZQaVTJbTRt01D9+Iv
nTlPRI2KKk3SXJ1RRsKB3wAn+VJDVzF2oKnw5IJHhIqfkJORKT+Z8sFNfijoZyuJQle+BzGEnbwd
bUOiCjrwBLmtKcPBthEhikXqE2UDKomh8bGjsBuWV4uUgO1qPMq84Emb4jkZY5lbzVawWnm3GOq+
6T5ArU4Z33FGA5b07inrWH+CL8v4H8/yncCrGUy6ad96wr/FAZumUGZtJKHj84ZeU3Z8MIw9Cvh1
YNT4Vrlm7ifUeBYCsOqFU7dkypgMkygxb1uKUg2WtSgFJmjG9vOZkfywzJK+1L+d9fzWJOTDvhc5
yOW00+XTdUMLk5vuCx0UnS671WSnpiKYh1/I3/oK3ZM3HAZuytc43ivT0taGY+NpPZt2lBHCJya6
E3mP+xV4gCBiZmbvwvotmy67idyNeyMaG9DLWA4DIqovKyIkOGlkZB1I/oCS0nsx/RUHAVGkfj79
P3NHNVPBaofkEQmLffK27MCGGEK0R6/Po0bGAzOr0NMhjjsxGhTseSp8JGC22zVr1dPdAfMNQoAQ
uykQcs0oxxuKxHSKuxqBAPf1nKyUY0Yjz78cSJKqJ2pkSfhCtb9AIOA/e8DeWjx84UJRBsvzRvuI
kvEu1XupaTleU9y5soKNa3gSYfhrfwdCpCHooG4Xi5WwRzV58MhJzDZDmIriIAb01SqVbbuctjqT
cywbLi65NP1ttdWygC20jzkzH330BgUUS1iW+G1ecr7+eEGE7PMvtW73yIMhFHwn0QewdYaZqnHR
81faiZTkbWDl0iX1mIetPd4jl3QBd1lT5N4YwDN28BwNtlJihrY7oXS+cp2pwvHn4Tqbir36oazO
4ffpELCLk+0B85GOMDB8jDrIxH0cXFOKF9xjIs+liCxevzMyMA1xtxuxzAUwtP79Lm7gz504od91
kEyAtwLOJ51qIztG88txI55nfEWcx4qrswAQJvjXgPW5F8ih2crgUnfpZ4oAG/e9+Wl7IRCwzeKc
jiihxT26pM+ihdU/pgR3dZS7ddGjycejKEs5uuLP9MjGC3YorMHRIGJe2HLdDEkjuyxpqiqksGIt
jT9bMgdpDHbCX9WPr9ffR0CgIhebwBNb/qD/Sia9z9uLhnkcZ1kJ2b5YiaSF8EG559h9w7ZzKsG9
DLPXjWnyG83jZUkvfvwo29vRWmTNfQ5BZeIoq5Ovk6BYVkQHI/LiLeiJNMO1xRXtIoA3l7iKvVxJ
GXfd+jy28ruojTAgnT+vDjaKPyuZXMML0RvntjwCEwF/mBCzHOsLVl7JC6NiH4Q4XiVyL3gkA7md
2gFhkivG/qHcfdU5qNX8PHdTUE0lhlakSaB+jW4LKTtas5AXqIaCsLceeTQ/mcXwD6k+61wjKlpv
uQ4tK3hZZv5nkhYh69dejbge4XxJ/qIbZUjYOcTSoTa8k1IIqBOqptGeKUVtRIkct0IZTj87qTxa
pbm7zLQwkPBg/IoPT9//CmgOW8bHS8DTMHZTW8fe9tKare2KkBUVq8GSoNT735vT9lsDLNir/rIl
+EDTteSBaO3iANk4dcrpCLF5pkgTZw1wLBoqNTJUcif8G6a/B+A0g33CMXgS5qSVQbmZegPihchM
Fxu6Pso26DZS3Mdno5lihgT/omXjLYsNBI6ptrbt8yNU+CGhOj1g03GcQzBe8ZPYJdk2yP25f4Ey
Ds1XFc2oK5UdPoLAp1wd+9G66Bxv+Jj21RXLPfB6t++2QUtqLm45WwXeeeFHZ33l+fGbqkq0jBp7
F/cYBGwfH9qd0oUlpZNrgsNSTY07e+e25MnBCWBAzLnpH8Rpa2wQJYfoo0th5glnF0/0MbBobTYF
IND9V0iWFt/XeAbLMeiwhLKpXPCyFWQ8RzNqJzEnSC0xBSo4749FPQbV2AZGsCF05l6msU9p6i6f
zin8fZzK/37cI/pcWU4hZ9T2r/z4vPbnh3/G8zNhP4qQ6nbIYTuuZSeix6qaIMVwc2OcynRC3Okp
foqz4/xuW7CybjqrwUwoOcCbrRVC2snLHfLCVs2HTCqlCjJ7rpeyLhs3r/WwfZ8vePbNyLIvEKya
ElgvCU5auMoEbUkzM9aw+E+XHSOM+nFnQpIsAC5MvsUAjBQOnt9l4naiv1yYxf6sqxaLmDLkDlR3
zZh4SUd+7maRRTXKriVIFN4AceMqGh4TjnL9JukTlz63f5KMkB1SOZveS76Si1yU20xeCjGtcOxR
barr8ooYWp04hMJOuxLtFKJ8t5hpfk5aaZlahxzgWI7VMHiQwE+MovKfZocDYoVPrn2xjEoeipKs
X+XPwr9wnlyCcK7F1goeT5MQv45RSg5tOLp2jHd3Ln0ReIgDhGs3261g6Tp5oy2MMgoKdjHaCVn5
bNqHaaL1/NIhl4rOhSGB4fjfNzuuZ6GtnyWiCd38Q4grZ1zv5NNwD/LsVH59HkJahoqxe+N58TQr
LyL9uOW5PHRQZsQxkn0ai2L6t1+GSeZ20yksmjgjejJtc6ydCwkclaEQGA9QPr4jsY8B6hANSbvC
z1/rNQn6+3DF9iPD7J9VfbwnJK5uZM+L35Qx76DDX7dqJTrFzhMYaqYuzxItQSLv17Mu5wJmM7K4
b/FBfmAevcZhvfIbDU8M4drIyPoXgR5KV3HtCbZqwPPkr1MEpROqBU1SD8mR9Hd2ia06HsSwttN+
At255/xO/0ALVwAf8OHACC21o8Ji5Jk4nQsLICd+jWsiVZlxZxDXk/SXfmjQCY38ZWOATsxtv/f6
uA1TxEKM20V/NqKtxeplIy1qHE5hBvdVmZ7K0ognd0iNH7lNKzF/KzEzfis3XzLpYBl2MVr2Y7a1
7e1SU8M5Y8hKaR3wR98eXpd+kvUGze2/GsrVfz4oen7PWWBzUc1nYHGBmrzjbExR8FCHr870E3th
iff9TWnnT4SH9T5diyR5hgqRtDKpm0yTPCNRYIXDWm13OgpzB0HqK13LdGNixcyTG9maR6Kdbw7k
S8qLmT4pCt6MaLjdoYAint/8W2Hxv1upV993HQw6HeKLA0uE/8KG7iRIEtehTf3pJkj2XS/hnJkS
qANh1K4iEQc7hQQiFKcbw43XDFmO02DLya312MS2nSBHGPwGOK8M366ZDa/q43J3lqtE/krVrlhJ
OZMhPh3QWyrS/r25Kx+D3QHmGNh4HFcpSvv8gT+yEquMwzwaSwcIXnLNNV3AbYoFbw/MU3BCLVDW
vSMrdxkZN3+jnuJc02ufgT2C4Cn5AlA2aOOTVUb39MWp+hXgP90bsAjp4pjyKldLZh8IGMzV8RHC
BGrkcywaLqFOFEGkFpJVZrf8JnA/x93NFCwmxjQXtOAGOaXtIHFDagMpxDAlNWY8Iw/UBiEf0td0
jEyBT0BX4tv26WorpXrnIV7BY9HUsOVm44sdbn2S3skTRPgaM1Gf55GeIdWX+oKgi1uu1ToDFO4E
j45JmdwjOxfTplks+zVe/TNmTaC7dKe6W8fCOfKlDDrH4TRauUwp7LMlv711BaHf94zAghysKgBL
ZxC9jFavXJaYuZoky4/kTexfST3wYAQ23A0+qtdx1IQ7KxsDe1BbCFrptHwZoMaKyYWMKejXTfzm
vo1tZI393RkbEQ3BqKgQPK5WInk5yMvNtcI9DEhsIHABJiZTi9nQ8aT7VMV8aGmzpsztfCYNdL4X
61kpqIrXCC66A9yzNUc604RrM2v7UEk2uakmyomg392fnpZJuG0OQ7NkKHSYlLtgOy1lWzCaq3Qk
xCL73boIcLi2B1TJa6x6i6xrzZTnPKS64fzpsuvSOjljR/srk7x6Q5Ll+mV+KqxrxFEYdN748h/M
eUD7aYRNziRxKi6uvbLMmTvoq8BsZ2BykQykCycxgkiQVxJ0Vv8a8LbazMJwUrjguVcm+rmXOadd
qXf0K3k4GssHvFZEy4A1MlFC76+0zz9H3r6LObQaAhQ7SOkHlYqI4tXCbtbsCnfgTOM2bFnkQSUh
9/0UdZ62r+CiA/5lzAffbWoAT7Eofqu6Iu/K0z4gR320elgSpfzLGp+yttNq7YcyGiEiYXPd5uYp
/uH45sw+snimgBFI3TcYMq3Q3xkMA8K+r+9lCD3cQwTZdwz1DGVwIv4bRvh4WiEAG/mlou53Mgcn
RHhVhcDlnpFhbazJsY7djDCjmmpuS78bYCUuYZzpjlY7q2XDW/BtLP1zSYaMKEG/5qfhrYvjQ1wR
fPSSyZ0PtyGCc68CPwsbCMOZpx8KYOiLMS8SJzoTAzIkJP598o7HIQY9DILNIz7C6SAdh8Qsxq2C
W1A2v6py4YflVTo+255RcokO9XNzsecu6VlwF1T82CSe9VEXiN4RWwQg3L8Z70yDx6UzzRIaPfmp
b+8UQ+K6t8lA7UE8hYHXhrDddzlxN24G6yCcE3JlqtXjhY+lZNk4KeDHLLmSH+XvWIzkmcaQcEar
f9qIka0rStwWJEak24qorSNKg0AGDLjE0oIQS0xXVttGpzmJ/WyBRDT7iL5n23XaSaZIqEfqiej8
mBqXUcf2D31dlpVwxbyaPe9iTIEF+jc6eZN5z1N4w0wdjOX/XwN5qvkpzX0MATxosML3JVs4xF0e
19kQ/2VgBj3Os8xzqaLkhGoB3jdUQaE/kFHjzowsCo0r2pqWgPz7N5M/Mi2K0ezXYnWIiLetl0ip
9ikimLkaYIUSlDLn7f4x11Fqt0fldBJbCr/7GaOkKNS3Waet4uFtSmPHcasy9C7fP/lqMmZVXCqi
o05Rcsmr2+0a0O7FXcusmPk42WyrUz+f2pQcPPOd0jK52hxUKUTo0uX3PVLv4Qfn/HBUcUVmgXmV
2wrBxJt8ekKU1okG3nNUlwc06lNhBOeSdibzdYI02BNpftgMTI+fCXg1aqkHoMLKmExoEBqUSyak
5Xfmsk8Krq0YX9i+X8dFWU2CLvT8iO4F9ualY3vg6SLwChlNo1fj3vX0Jt2fi4uusjFSHdHP/zUv
0Cqk21zjIW4KlTgxsytXds4IF7S0dWCYQHhM5pFxHqfcRicuhC8YCkxNA/+R5WYVHhyk/ZLamMja
J6r2oMmmr8r3gLaTSceHmoFyknzH6Ld6ncpmbDtWo9cJotBzsvCwmPK6KOmXKfLApn9Qros60Wf3
PBN0Z7jFOBP9fmXzplFqDJMjq9Uft7XW6ba0fqnF2z2zvFHi4Bz8I6Djj0WZ00xJp8/EBh/h6ZAC
EQZI9qHGe13Xe6uOzmxqDT99CtkLtxPsTeHy2t1r/v3cSo747UnMX/ec4Euq6UH7hPHOFKLY8Ffq
xWkSrkbwiLKZZAyrrfftIY8lYbI/+gcHzXbalgP6ox/nbUqU5r0sxSfcBkk+fnt+nvY2MjHT2l40
9yJz8uZSG+9Hu81NqFc9N7+ST+v4M0JrKorxI+KaXEnjEIIH3fpkdgtrcBLNJLZ2YHKr1F6eGXbZ
CjgaWCE+dotSrYW2abv3jXgjzxsy8YMX6qEENlvxIPyrAvjtZW7GXrdbtqjlaHxP4h5RQeb+Ttq0
vu2D0FYa/87nhF0WsLGfHMGa6ztrQDbvbDEz3imK4jmdNAQnq1RuO33wIqx9z6CbQvqyfg47muff
HDIWCCaJAkDGm62bY1gAAgVbJnVmhkkQ8y4gg1iyFIaRcCBZ/CwwO38MLEFi/6TCIImV/WEHhVpn
k/17BJededWtcFsGXq+dhK2YBi/Y6QL6WtMbREk1Ao+G/Uekcu4iw4DUCbmyHp6wYYIFT8VM5UXL
CqMV8+dk9oRu/a4vRHoXG7oeOcxi7hLUjUT9Jvc5EAYYXLq7pX1R3OFXkl8gXfEY61bA5b7r0kxS
J6WHjfbP4tOGI6z8tNEOdHoaN+s9mdkXd3glIQM7IpmQgnEE7L/EEwVpYdx/pMuqYNTTC2gBKwvS
FcD8joawABbOx/qyT6A3Bz5SYOkTdVr2YYYJu2aFrb7FAdFzbrb4IiWaMi9LgSIm46fx2k9WLkol
3tYhgJuOo6XK3MRUir0Fl2IASJMfNxO4ZWaZwFUKBNjZqZ+8I/9rAyzVrph0z4kVyR+fc0jSNvX2
Jb/oRGh1IXh14lLjIo6OOU/X+k3kcrg9WXoGUsozu02+7YxfjdPYwl06RI84nfLQl3wCIOTCUrV5
qi07hiXO/YFLx8oiBUsp2tjNJkLjGlwqIl6Xs/TrP+BkFAGMi7XK1SaUm74opWXOqnOrBSx+rAZs
BlWxBz7gByiLmHFf4QgqBR8/qhcrJrXcvomAdgZW2tI7OhZTBNqzZODtyg8rbZVpicoR7KUDB5Nn
gH+yX3RwzwUOAE6MFSs3xgOa+5a2HU1ML+b+D0v6KULA4cNZJeHexPyWJvJzfR0qX7g+upb0r4xZ
isbznGCeaQhuw2VM+NkhE8QOjTmdGolUwfssiPBFK9euCd7d320mgmEAdTcAxG69xEgmfp4b8hae
1G3ou4iIZfiabbC/vitITtDz89nAUxM6roDfb8KV8+H9y9z+ExDdEqShmfg0pJb9Ipqbjl1i/XNI
hrQgzjKEXyuKhxe0y+IJfY5cr8MtddrYPUKFnLGYmH2uKAUYXbtViD97tSMX8tjFmabb8xjNHiBw
6L2/MszHoonCj3vToFSso0qTnX76VFqLnDyzhsjxnJG5NIMxOv31ucwjitFWWrphVc42w2GiNMoS
GD3zmXrBLsHl8Pb819aU0cB6zyI7jYzLb4wtK98wl9ovjB8vVKBb9VUnN4EZvThe5uCyoNC9dq5o
JrLKHQqYF5EtNwgIGsSBUkFWfEqfcVu9KBWliDzi9RpqfVZQK+LNmoSbkmP+MUddMd8hYrGIjxBa
F2qtLF/kXZl4GwvwJBpU6Nul6CIXf669xXmeJ9tjCfkE+JssUPQ8HO9nqeMaUzJgg5nyG4Kl4J/O
drkyvhiWPprz1pw3RZn7k7LpUqINovBwJUs4tBpWAAMqgMAWRC7zK6ymZmX6D6PcEfe9LX1kuK4D
zxNlMjCFLQRPk0VSX1wyQMZiBR2AmNmNevGwrtJ9DOEzwCgPjKGv7nJzC0bVGvFTNf+3knX3dA7+
0HOHqlr2r2jONAWYRGCWp9pA5z9Zlx9CNOfgPC3rZd9h36UTTNIQvGE6AY1MsYPD85+XfnyHh3AE
dWu8U6uDqOtZ9qyO3B2HoPFH/hsjrJA8h/l/bE1q5+p5jSi5uPpFRnEiIjWwpC3y6ftI1vnvB46n
wdAYAp6v9lYigpFgM0/E0J0R+HrFMmevQwdvzaIhwbWSbRtQQGP3Jd+M22n70HZNyuhiTmvuq2q/
fhkoB0jXzX3tom19WanKOp0JROuTZZKTCt3GaSZZdTmgF1E1gPt0i3lx2Iz+NLlJV9Amb3PmDORw
2/HmQ86UWE/Lrn9ehkrnAEsXy+o//SXMp91vR/CGpT3UjxapgAvjZ6woZ01McKLye0vKKD/5WmXD
mx/wCmBfa41N7bwjn8mWxL9vUwhaLjhKbDfPRz+mkMkXHQJZmNuUa2fVtlC5m9KQtP5947rQmkMj
J3+rq+dLY2x31NfjgttX/6dZVMPB+JCcSnuzCTK+g9GgWHS5R21jCyrXQMFw/q/nTtzOBbcbCDx0
axFgFKTr169WSNXlAolfyD4xtCvmAKIHNKFJ+m63lAbsuld319DP7hNyAl5iAnkCY+UzIz2Vsj24
qvZ0ph9vT9of1aSaDfYcC2EYyBe5HLRq2phMNZe7gNnFSDLOc6g0CgltJ/e2HGTYS9zR/BXrsjMb
SDtBjsF1suJvDIDWAJo8lxSemFqYi8Uqq30wlWGo7EnvJQqOOUK/RpPjp/gQLaMr3vBqiPpNt0Fs
2l2mkX4/BSHFXTmnKf39Y7yI0L4EJdfaNSjKtJHlylokwGGA/ak3csEhEA5mJSHAIQqxXvrY7ApN
v2LJppNCRVtKPuk+pa+DoYQR555jVQNdzziI/EkD9DEJPxKFID5AHDdFz5bl/vbjwAugZ8SBFTRY
WvLhId/uNkfDCx8/7dV3+03dMjyPO9MBNLZEqbYzVCcvDwhT6AX67ik37K3kKRrvdlzreMzXUPee
yPefoPJBZeMUJ01nyrqDeGPBMaicKCJLtSS+dNEPEVu/thjCqceDmT1HS+pxKsfWsaLqewnBr8/I
vGulaV39joFDE11iG6jUggyuK7R9aqNnfMV6Vv9brjIbMFZaefxp2nSRtNq/hviZTcoy5GPT/AS8
3GyoOo8m0eBW1vRbmGoaOY82SIzGd2iK6fs80CrqMGGTacXs593exFKJAeI5TzB7e4jlVphLBpun
YA+zcgYid5P3S0iKRazCNwHbAs6t6DyQPkV9/3jd1VoNrDA8SQQm4dZJMKBm/9REqDWNfotC1O4n
vWlfscC2rFlEU/aigtdQe8FxcTaNxbgnZ8YwF4ZMzHiUjLnWaXXvdUK40l+vjrDKj+ezy/4Cbskp
0GJZHvqQG0raOZv1yABwo/PJa2WW3Y9d/RAh8US5WO7KCc01rj4DVnr3NiPtKHxrBKZvEz2+yx9f
SH+Nqa2ONFZIjZYqTkG5Fvyw1EieqqU6p1DShDnNP/XB1GfAHk7Z+BpKVaoSBjZrL3kUjCDZpTeT
N4A2nU34BwGwVkqNKSvjL8O9UUaooNx7qUfHbJ6Uc4C8go6YCsaAtPGmOGo6v6Am1fKOCJhxU+k1
1IYeQldmHuuY5N7OFf/IGbIlpJ0HWLrgt/p9FgNpQcV4ohXTHXs/OsfUBLfrj5MEsCN/Sd0PvF41
112UKM8AoTKVVg0NIQ8bm9FF2Ds6gFL1i+4sma6F6mlY2G1dtnzCZM1MuXrDfVmVlbFgxOEbapbJ
8UDrq96HG7agE0jCn0VIMvbGl4DmUMjWipvH7AQYJ7u6XR9+agWJQqnWl6LhAydHmdQUzmvpIWO7
x6uCiO/d2tOXnVPrNJS53phCG9JwnBx+fDeDVtpCiySBzk1GRb2/94ZOg/ZxQ1l3grzbmTPEOtEU
VHw5m7vqSI+ho7mSej6az7/WfeESZdmsQKj5Mf7+05X8GTlYenfFVaZkqoflvcqyIRGg80Lls0x1
R1oNnj/bzP6fZMVv98bGvN5/ezX47s8aVssXwUkulPocDWFjE0JvUtkMYx+eWC2TGpy7uaPWy1dw
tjm6ta9Fuvf6mCyHA8BAP0BlmKzwGpcWDFjGqj/oWnNBjbQvtozZcg50gKOulUsCUMwBifMf5cQ0
AHHMEKXw16PTeC3fbFRstujqBBQeBeZYbLY3e2rzK6z/bQNAj657zSs5upNwuVxaW757OsokRvvL
f6ae3v7CvtSIuNL12AVD0uXvesSR2rm6F0KV8mAw5KzYppsahmkG5zeMCnRRldO5gMUZC7+E20fg
0zRNhLE2ztsvZMSvVG21f433M7MeQHkS0sgMOIrqP4Bu8c06vo00vJepkxUpjOuzCvRoEMcyXZrG
8h+CYGCW7TvCsVudD2AlxszgGrh2YGTrjkm8ouPhyjtxMuclBrj2Jo6y9UUrAeMTPdNiwmDLM6Kv
EO0JpdXdoATNA94y+L9WvzLj+XX1OwBiie9YDrIs/s2qM7rVjvTvKt59Hw7mwre0UeUOTB4mX0w2
1ecEt5/xsqXEprH7MgRYzMPSgngslZ4OGYfTuBREQrMQzkVmWOovRmfiLstEVztQriiKvfhXjqLi
ZgdDV8zMBoFztApo3gAM6mmnM49YQNgxE6SDhtsFddLibL89b+ODCsG2jjTu1aVUvtxUOUwifq4R
6+fAUteMz1FqEAdidrrC09lDM8b4BknftHvTIGaX+uqEZWClzpHnjuc2Nhpn2F0vkV6yrVQoW0DN
xbaXk5I0HtK+isrX+mtGk0hXIWv70lcp3GfxY0EVmgCJ7l6i9C5ODhWRfTBB4AaB/tE6ISXe9HXb
1f1H3tYmf5AAc9ZmNizGhMA8McGELY53wL4N15T0eloaPjhRvvoBiZlV28YZJP/khv2lKAEbbDyY
FDtexngtxrEaydiPvb/RsiGwAs9vBQg2Iz/f0Jgp0FSzpQJFgFqmEArLHix0ANthxB4DGqEbbvum
3wKTe2mTxlizqPcgDrltqIa9eXPyQiLfSOQW8OAYJ2shEW4zxKUPQHvbFgUxakevJvDsNKQ48C4K
Xa5Gq0Ti7v4svDBicrgccgQq8bhfD+iN3TWrXGQRxKzbAshd86VmGBguadL3BwH5/r/zOjZSrXHm
iBpNE8+s5ojPOW87ryWPi2TNmtSkkyFymFB4j3KNdniSzxUizqWIeAlXBX6oSPBtOEgNB8eHLLas
2bHsV3sDQFVyTb8go/BBzHmq9gi+BUQAgIN3hZOfL5cfACUDyOYeuXxs1QAwKl9ZFhys9+9BiO2o
YviDzqc3qQ8JetFSdFkHMQLsyUxIPeDtJwNozFY/7HPBOWTPkozBSmk8h+gfEJMXpqz4LKoTC1tD
aYn7BlXznMd06VANsMyLeaZ7imxQLai+Vu5FZ8Kmf32JOPvMSwCmNxEzXPzGm8izmqOu43f5U6tS
TtjOF6FIayQ1rqKygI9K1u5D78loHwLY7YvxGlxfeJSGZWpQkOBbpbw4F2W/lB8obHpn64Huv+zb
DTqCqLdOxVU5T8lnNe2tanmXbJo7bQPQdYa5l84ofhcSGLMlvY/Nf21G8HeiWpM811hhwpdNqfdG
A4qZG1ubp8LdC+NAH4YV3KA17fVPoWxQNQtnmUWQUHCd0WgxJXexIvQnubvRgGMy0yjTglG2whWl
Utby6qSxKO/NluyqtoBnnArTUmhNq02wnFwBI00nHsHEQ6DYJ59Q2/7WX3s5xCNPvQP1UjJl+x4O
BGu2/yUcxxi5ha3MG4lUMLX0Vk+aiUfpl5tivgaHedvlU5Ok8hq8Qb+6oLjBh7NXJu4uD+5Yql2N
8XS67YQRuYa9Jngqv69ZUqNaGFveavahXIpUB9ePjlNlWeNYVMV4168WYQ6wAISJ/+uDSeMgrPtG
OrWxH5jpq9+GyFqglYHwB0GWU3bI2owOSpb2Yi5X+A6jBfgl2kVqLNf430sh+jZnmCSI05Attn4+
7Vq7hSFAtcOV3RlPgVX4HbuUucNrCSonqf76IwertXY1kgPr9ADKphoLJRdvcTDGpQsB/ZWkCoJA
PgkEwyr+rQR00PCdmM0Hx3qyNb/8pa2is2NEqIav2gpUQno2KLUMLz2+dxfeZKrnwVGOBon1t+wp
EeAeDH+h55Y/HsnhrmBXlc4ANbJ3yDs5QjZghEw3Ik/dqnlRI/5gt6nMv+s6AtsGfQUxhE7IXBy0
V0g3iuMrdEL3laOJBjCiQDksAXHqUpHCN6XwWiMWp5FCntIdv2aI9QX/SuwSIheeWt4Loj5IcIQg
fQgvCiW4BByVSD4swz5hDr3TXyAQmXbWNAko1V0fpIWhuGA9Xeyx3at0JO8vhBei55YOOg8WEjwz
r3iLk9NXzeSK2TpjKGF3UBA2MnrLewE8dRpw+22iJpbVNnPKB8wYzweOCMR/xc2l6QmMShoxDpXH
BBkyhj1z06xroz/mGdgd7Jszad1ak+CtEacvACDbiNWF43GDkna+NJWUvKtHpiNOGShsybkGB6z+
AbeZh9b7R5spAyZSXmTnd6Sl4VESM52Pg3Qqa9uCbvpVfdaQscHfL4EcGyHfRrPjZVKRYuPcidG2
RPzHFZH+b46zdg5+fkSwvIDEGnrFpQ3KnptRT7dLqnmTcB+e7ifOtMD0jYZDEApDzi11dzcnHaN2
T+ICB/tvrHdV9ODkPNSR41IRe9v555FucWbM0NnqVi2UZZFKIJh64tN0Q8tiWddyzhZCmWgg7Esz
N3aOX5Ay/BE2d0aegHEAbFGobcnIlcCuntGitpXJ4dQHR+x/r1PX47VJrj+rQR58j8l1e4QHcjJY
jL3Vumu3FB+72+6GyZOSarLpfmfYaq9vhMq05nMQQ540UJvh/NbHPSxJJK+Z6qtbiID5F5jOZRYV
ntKmhgqKZx64nuQIgULdFP2Ssy6wit8B2fjTNSpfua/3YAOFD1KeU/1wpIObIUJmpuDE39XqO71t
2gQdoDIXIPRzXCc+P4AtFd8LSEFChZTFHqt2Mj+bEB8nIwYzYggfczZ2Lic6rNzarRmfQyPNvCKt
y8larIKm6AxxwUIt6Ojon6+JdEX9+VPXRwqUVJNYYz9mwcx/pSbI1VUd5k7ncmHp7iaub4Tv56xC
szbeK6PrOb1ToBJ2nmG5KWGtkh27IHqwGLzT/GhqN6PmoenA+BL8BEzwvMshOJqRcj9YqZ7TYflK
Zu1Gwx93lZV8UfRK8kKjvCfFSNdul2jMUd3DZ/OPeG+i3zAMoiEwvd7d3G0AOXY13b8ovEWXZUjX
52UtjYSAqJh6il/0q9FwL0hFnS/DyNsdH90RefeZgFZyy5npqVtXo80A+Q98DT8kO3+f5g5wvuZd
5BPFCq6Ry0zgNJZL9pcrJ8T0Ab4ngWrelY0/XobZb++IVE6WOIJvA6TihZdmzzQm7QSQQNYeT80X
uCgylFUxop7HyhQSU+xFk8ge1ICAZvrLjEsk69XYBrt6ZN/YdRbIMkuPHvA7q+0R9ahEK13tnyAz
59TikH/MH3kDGSVzXBZtsnGwq880kk1Nu/QH85OR/u6fWzby90Q725SifDPthY+J/W9wJXfAPYTu
GwePzr8+XzTGFklKSkd9I3tNGWhaaNw9WYjxOEPIPlRjBgERnOMw+uCcSCgpc98hUPHKAlZI93Y3
sLNyGFjHc7pklLEjKUbqhunNPJcMsZpUdP6EBYg4COEkfSW5z+WlCKnGUDKxFqAh7FMakxCi6s4I
QzcM6DnAoTMsPoGcZ5kZ49Xo/9jF8WNDrhEEkL0i4QcLuwPoiZY3EH9cZ+VwSlWUR4VK1XO0sKlu
oyKQRRhzY5pmcHm+saeXL2bWAbNd+lYbQwDpnKAPR5N4tuAXihr+Keu+68q9tNhQFKfgQZJN9UiD
xLpaRTwuIegrCf2ZP35gMi+ZpRmt3OjAecSgvahnup/l4hFVcowR9Xecq1PcbXSLvFP0zTBlMjrE
9wjgr9Pkdk2bp8uWyAESCUp3NJWMNMEBnPaGXR9r/fpqnfuo31sQoZ5nCu4do8SMx4mb/mNeEtm/
aX8HJ/Yyy1DhlaPPTxWXKzhAXkm/QRpzZN662pEFwR3JVrLZ9AljXdjNl/3hoAV8SYJbgE5o1Gq4
d3WkxZs4Ypp+KBO//4OGoVFtAr5Uz8jzCAVeXnZuZu1Mw5j5iLW/GubsA/xbVoy8fyld2b9CN0zf
juAhmnLOGyZw4JsxPR5GwGXBUnPwzqLkqngBTq8JJe8aM0y2F9klB01JzESOU4kj2hU/UT76+Ug6
7xP4cqZ9/ZWu4/WrL1rT4i6t7HHE9PiY0WbkXDkEJccFIC00A0JzTt4N1K4wnPqx1SSJSQ0HA8mv
vlBF+79m+eYTRZUj7tIELm51MEgrpAY+s4/pbwsBLAaJzbXeCAbNamSf5wkRSmoDO6ismnuhMtup
KEmjkevPU0hB1W7VOcKTA6adtTZgFpoImCsUIewTit2T0nWlfj7dsKoKRGcSKxc0YcUWpc0hj9xV
qdElVwJMM7WR1McjZiJjEQN9lC8IkXRW/TrAOu7dRAdDoA6bjRetrMGlWZNLycXZcG5N8MbU4aPj
6i8g0Dat755LJNoRCOlBNFK/LpmH16MmkbDcCas4QajNpOtXRpL2o78v5ERm41cLdWkxMcncq+ue
lB0FB7PN23a2/OPljnJq9mJU0hmtIcYwhNwc3jN4Q0RgRwZZwSXblkRCrTPiZwKiTMNlD9Tu+Xkj
tiaToCyYZEJmngYDtRsZLtJ6vj2a3Olg0/pRHXe6QKGZ2naxteDnXxFQHGOSy7qD8guq81AYoKhz
Yca2+Umq4hmmx5TBMeZ1HIjw8hC0R3BHjjjfMXtUjafWCgUTUmqu+AU0Ep1KHkVoLCo6OzgE9EnH
tZT0oCITKSZra09zBERnRXq2cuLIxymItpUhiaV19qYcaaCqbE6ivqhybSM2atCog+sK709VyG8u
5UqD55zPPpVYihceXXbYjcqUCZHxHlPkefO4bp706nScTT3djSeAzmW66/EtCAcZpQ18ssWCH+QX
Tp6zBO/n5fauBqnu+FJw+2wElrFvBr+TRGFfIl8JtjpM/i9DVINBFsZYvXK93EY5RJvEHga6t+93
Dznicy9EFrR475/hVUORzGNVnpiHRgx/BvqHczKqZN8CScStwjYKcFbiPwvc+bKw6sWIT4rCHR5K
xY6LP/AGGAQxTPBAvrPoSp3hjNbkBET+lj7CM1gBdm+/WnlXQn8nvEgq9G151KUTV7xYAXDev+cX
MN+oAa6zDbOv+aOzmUqvTTYxZv86TJsNB12x5au6DC8plV87lcqjJ7en8RJjYybGCP6r8SZkKMDI
B6573PvE1vl35DuTD+larTlrQBx26K/yJYe9OHZeRrVeAA7o7YFvuKtu5OxtUT6lRkBuYPh4Sx1x
UXuw43jlNVZ8G1cozyPLKoxyeCJ5M+FCHtcs9uRB6c8vEP0v7PbE2G2jZZtGhMiELnrjP+1MdA+g
fIZ96xVwFlMwF3HdhAtx2klQuGPT1tuDgOHKaAsY2oyx370sbyyoULqsCKiS6LnMYRq6j0f6j/rS
BMVNbN61HJPS/FGKQifVZOA9KavppQTVEX0fPejMRb8nuklg/TorIaS5hJbeFPHau556sztC68lX
4zfcktjx0bIcsmmXcNKqkEuiLjUUGpTblEFl2UmDe3cxvKQbFpr/G6ZetH7iF4wwRHlcAxDKFUBt
29cs8vt8Pd848z2TBvMQE3uUY2zZ0Ys6Xfo0AtFWUSZRN8Bzr8JM/1F6dvuPOqf1qXVN7exOpAZ+
Jm3tFrKB7JfF/VXWX/Gw4P1W7z0iyh/WaxygMzMH8lRo1YbDxprgj7G+o2zrToj2zJeiruXlnwqm
xzLkDPzKuHRMhOfQXejJLSNnJWzgX6aAJNuFmBgsVRacfjFjsv4zIzoD+LV8ynPFUvryFUefx4Do
Ma2nVhPWWILCNBayHSob4PglWCFqb/tPQl1yJKb1uNm7Ni4LIjOCS3OIkIVUd3OcSP3LA8tDNuxT
NfyqaEC/MFol82xDfIsssPa0LcoE4koQKc0TqAPRaOTpFKKmg1GgY+OAonHzKlN6XA51fn+4mLY5
AqtpB9Da9bnMzqgB5gD6jGSAtgNGcb6jOCHDcL5gBrvJK70atU9jJMAEWo1hUsZ04RIbWkNAAYme
QureSCcnaADvfqDz9Xx6SZTIVXWt2OvcSPMvaAn5erVtHNjTuS74E+GouPnw8X/uj5pPT4h3+Ln6
Y6psp5oS4qo0P7vcTncJ+YlG/OsfCJk/v5iQKLS+FydmDn+WxXGpV0ohrCsWoV4sPHTBDyHuJC0W
6c4PORqLYaZh0CY3+ZztIFRuxkxAyt02dY1oWE3NH9/jOQ/RCw6D4Hyg33iNCHaHyKEbV3P01GKw
9dNy59835Zpk+45dcgvYUFTjZ4hMjhfTMoWts0NZncJNtO+zn14x1+rHCOL5k7SitVx14WZVGiGy
AAk5EGstd0V/AfBK+p0vMu1Kj4QXSNGTBB6qS8gu0y+qbnd3ViRXTNl6vpyCId7AXZDW1F+esdr7
sRnyi8Q5KqVHDKEzVGhc9zkZjHGsUYsibk9Rvpel/9kCqjPSTLKrX0qcG7u73sZFxngCxJ3HV94Y
Zr94B31oil9/kWoORonsv3IS/+jWdGaMrPJHAhTb1QFuejPCZYX38X57RkOjYS+kj+AyhA+0CmSP
5u92i/xL2Ak79NpHbys9nXYL6flPveSnrHE6Wkfc8WJh//USCPT9KrkespB6/J1S3uXeO81b/pl9
JChtUiubI5Xmgvtj2f1u0mswe8YA309HJDw22rXwX3z1ZzOd3AnZ1GSulB07z58u2v0W3gUhOe10
pNBZEE61WZny777MyNvQpLeGjnCsm3I0c6xHLqI+V7uNtxamYDQFWROIJCp4l/Ef1Tkq1KinNIyf
m4rpPJrZUIfQmnOqEQ6hjuzltpQDRtDEEJirji64ojTJoDrUlio0C9gnOu1LwoEfixU4lPnl//46
1vv1qoY6wCznefidqlF6cMcEVHisTkJ7fAz9bw8R4aZq6/nfx3KhKSRSlLMceQowAmiemYeqxaJ1
Uxg8BSnMpTNH5NQZgRIbirXvziBzAmk4s3dNyBoRMshzHeq4yrnRdjW19fjDuV38thp4kdIyUPKq
DaSn9Y86EnZA03ZeeCrVNyVIuZCXZrrA+808ydbSY/9SMbAZzMdsL3KfUNcZWZC45GPNl6poUJP4
MpOLBOTWNfU3Csb0yxyZ0eEviUwULjl3Tv4gFo0sPbKNWF6WfWGKGRHEDUC5CxsrO07iWmCOHhc0
s5UZktawB2iqpynOr1a7SZerUP13MA45Enwv30LiovmEgOQbSMWckyrhnTsgMqnkNybSJhiY9/Wp
rgkmq2YRu8/R8T+SX9Mev0ami8T/RVx4xp/yaIqlDp1R2KUPZE6AfHYsurhE/60/7vcQUazEUpEw
dJux2rFlGUMOUT6MpGg5mHi1HexXveoBsb0MPPXr/Bcn3chrV8BcoOmM4E6AbswhYqF/2WVwO3rM
I7OGacrpgsV/q6UkJDh4I1pR3aX5BX7YEzBgIlJq6bt8Iro3owhQLe5+YyEZk25o8XdHXT7UMiUA
WEBtXpiRAYE2YD23cCnx/U9P5/sG1uEN6RlB+EniI4DqtB53J2CKEQ101Uu+pOUS1HLUt7aCpAXd
TLUvsPC9NIUXgSqBLIMGsii9IDuHLA5+BvduOLEqGbhejSVONeg6AwFfFVs8bQtHlQTTp4lPRMWy
f582gzaF/jAWd9dwG73l1YtzOhEbMjlHAOlaYQsNd5Duh1Pg2977QeqoP+0J54MeNihKUOdNjNXb
/KgtrtlJe513fKXh8a/TA8epbPEwrNl2pmn/c/gakJ9Yhje3fRYgLPGO1Y2/4CopxMxNrqFmWvqC
LYksLsZquGarlVlG7uOGr6AfnZzfxXQgh8pu2jH4MG6EivK5ooB8/P1MYkIiIpN9Cs4Jyq9JDMuy
+2pHtsWVQ9UYPicdq2F6e/Wntc7pqxJnI25csPjPuv5cc3UgkuObEdang1P1ecnNiiJ4hST9dsUn
FOjvjmIcX7binNocowsFQ5N+aSrhVfOBWQempAzDQ6cmGao/qqrnzK9T1o/Q7vEgEa8X7oTrH0Jj
ue0/aGoc1my8c6jsSeXsKlz1/OSDdrbbd1c4I/EsM5fjXJRpSnfDA9Fgp+QorCAMyzbWXNbRN2QT
6w2g7KuFOana6jbMgBRiB9BKrM9P/dwS+O7b9LfV+oaD4Qbrk5Y7KU753yBevX/Oxgn2g0QBmxTq
gOdDKbThsZFGQjQnrFp0YUDHIDvDqkEXpS/PalG5SJQtI9ig5nS4DDCc11KT0xiYq06JltVuuyWb
baZggEpOBDaf3GbHR1MuStfZQHBOmEi/djmehlw846oQ9DF2tlZir+bo6O0WF04aUGYLsnK5MEjE
FDqwY9yVLZh6tL1id008JYSyTgZAqCwEHHWmOtbmtBG6Fv1VAk8zKStsrvfvdKuLG187HLoTXFub
q/USaEHoRtsg3AYzf9iL7ALJAiwm1t2AKpl08qyxv4NtRqsxJZuv045JwfhQ2FHKQB4SJGenUkTZ
0uKbhZOscEXO+CLgs9MsMcpT8dDd2ErdeE1poDfyJiULM23m9SAz0KiQCAADLWPprQHVDJ8LnK8K
qY8LKZfGS2L3eg4CEHi8qb6KaodnfozpMmXKtko7qHvkNf9mh35gJOekvWsIIrqkeVczzYfrGRJf
x0m4whOTQlckvlaLv1qutk+2m21GUvUkzBXl34qTduPaQRpT6YiPGb68JhywYqGP5bTuEivjecGF
IFAz2Yg2Dg1/aMuw5WQ2D6FWfF2C4YbiD+KM4pSAG2c3i9K3Tk+MXoXLfjh8tqC7ckWWqNJoKsfX
dJRF/U/ae4FrEFVNVXiOQy+7UiSqZxgDtGWIL8PYZ5xjFLPBF4YDp7DI6hLveuPQKV1ZEjG0P/5X
pCEtnYIq41x9csOmkt3gVmVyR1rnmoOeSX0s7Ynh62ViSM+9cW3CAEm+YTOfn5qd377JMFruqCK7
1oz0caKDxMoKOBuSFiVBxT7MbOoV5GtSwVPO3UBcJQg70jjZkaRFG3g9gdTFDoPr76DIVvpDLIHd
mrv5086Rf2o70T5bOFcgHXcSUXMii0Cqe4SF2Bt9ECmMxLMyPlb6MrfkEFHhhCgJCS64MD6uWCll
O5ezm+p/JuIHZLPoStJH1wA/oY2KjTWpuZFd4UDx931Y+kb8+xc2gmLJ+w0l1MldU2mVUg2DZBuP
cz6nu0KqpXJp0Fvz/Se6W/ng6WDOhdMC65e5Kjf5U3T7VjXlkiEq67oTK9zopZn/RZlxJIMQRPwN
Hir7Vn78UxBvJPM9DdHjRvT8Dx9Ay2/4OKtLkRp55g5LXDvDNm1S+fpgBnGPfJdyVBHx+jOmP0ey
NI2La8AHn17Xy30PyOZjxdEatLikhRgiLhIMupzIwQ+JZm/dK3DESYgX8vUy+FfXcIf19TRMrzkO
X+HIQCh2K8Pcd6+ph4kEUcQnWencJKNNTwGghwOqsNc8a76yNIN3kX+AB+k8ezlU2PA/qVRhFAgO
1fM+0aPpoSRZh5kI/pZO+yHHAZSXzbb1lP1KEh2CJjQkXfSQSQ9dCws4SwgbFS6tfMHWNGERL+yf
usKUFdr3YJwm9d2lyAqrTr4HfinFaNpaIjGKY/fMSUYesRrLDB//bcwx+5Ry+dwH8UO2E0BPMwss
0iNbbXTaQxHo7qSUDuQjHm6WudJi73acHGKrnj3t8lLp+qzXjxWgiu3RDwtzKx/OAymJfhY1YWuC
1jjOw0A4krpwbnvi+AHthBoHi0WoB5HNnBw2zG6YwIo2S2oNEb1GMWBf3Lf7Y3oDoMOTKDgsYlJw
sx+enEtTCZkB60rjC+1B+A78VfHx/SY0cNJiC7x8bagFyDxEqGKDyUpJSyhvOh+5FYlPeBD/5wRY
cfO9CyL32G8bjUss1m5DqG6kTP1fQ7R32LmoN7Mg+E0nBr01rEdjbcMsK1IaGFjyoNqjA6P2RnbN
FnNM8MHEQN+/VSFeO8KIqn7WONQ0nE84L5CGJESEpos+xOOb5/K/FAp3Rq9XGVQKXrIA9aecrxU8
zLbC3cElAQ5eqe1yQy1NfGJopXrg31F43fPFd2O00W2DkzOAPrdEShItkHFddNckSCsls2NATRcm
5pNm2OgPQb20YH5s7lRwtXCy53hmwvDulq2WGfnE5V1dgi7fJ5OeeZpKATbJCpxKvRT4/kmx0gSE
2J6HtHzMni2O/lGQUXP/m2dTeZ9adIAvG/KsLyGK1e4r1Sghk+AlFdR5mYwrrXy+pSaxfHaYDraf
uLutBlnXKaKUOuzbmMV2Jnax0TC7IgJ58vdKoU3TceJqPNUG/p3b4tPpfviqpx9psZcBOCXFDQjz
pG2qj8ZjLkP2hIP0mZygiPcJpwi5YN8zLWeSTGoaQh47q1qc220PpasxS0oYsQQNw0vroIVPBvZv
ZRQapMK+eEktcZtNuii2cHEuhEly60Ja9/2Xk3IccKF/ETSNegYJy+ThoKRteGnIGYRR2KFpNKCC
3aMxa2VuYFWY1xTD9Xsx1pysLJLIvV1oodCOXXs3GSk4fHBV6MYeulC15BKeZXs5TT9cLz2u1qdm
7PYC+qro8+gJp/VSAfc2XzEUNOMwRoCEvAC4fINAfiR/FDxktekW9Krxk8GHX86yBubGK4Ca19Aa
D0BZMDUOqnEM4H88idUifNYggaKl/cdrBaiarDoEq4W5fvICnQH7kGocvGrt7L1ksFNfcze0F+bK
akPyBZFk+8db1LGRvQd6kYUHdDacxXcmjqipwfQtt+6OJ+/li7GYvIMs6PwRC8sEuABe5BQTvD3l
lQ6rz+JYjKnZiH2rCRwJwMwHuBtlYeSWorAAsscf55wWRlK2F2ATQTLWH7yA6M3P6/5oDAz/eMKA
P5HlOomJ1oeY0BMOzSSo2F4bxps7qJiMa50riUe0NzTg6v4+mBWEDxw9yDWZ/teCtah0xiaxMitk
Lt0NwTwifGu6h6u6NsIBx0qS6FSJRUAJFGIvm7Go1GJAbcIqsVHMGw1AOcBFj9cQaCpnuDnY/DDF
ri7FE6Kf4bJPQdKsH+PCD4LXZp+/mEoaXsoM38IkcpBhGY3hTxEvzmLuHQ7vr/Yr7yiM1yvJ7uuw
q60XVbQ4/iqf2HYc5PqpoiKaFGT+B8Gbu2xxWL1KBMRskCK8+KBZZ/ldMz9erlxYLDz2j17bUdwl
bXId8F0nHj0lafo/fQL5rQuzWOtu3TyCBNvh6teM9D7aRJ/V5zbn1keUBcCepi6dsvyaaV1p5Tw+
xjJ00xtzwN+rkxEI4zkCwLV2vufT/FcbqJnBewBdnb53GpOaoYzx8jyPz0JWIOeSohBvC+2HA/+b
ELIc2rjmeL22QtPOIe0pO7lPdbGieLqJVlEFXhY9pG6G19+lnVp1e3KB2q4/xO0i5BDC9Ce+T1OJ
nx8TIRP8A+eCoHkItV+hBz/UbfF9JH9qS5LSSkjgIBV60TAVMOxuxpE9NsA0Jht0C7ilZsSIaXYY
wptsZuD7fwwSpM6eTyR3QctpNa769ZvmywnQwKRVwsRg5D+/VIPEU1vbTxUHR6AnzLUoLmU9qq8s
bL5Cp0Ly6F6jtTpoQZKAKLORSI0nAJRRVIPfme6QzsiXuDqsfY5LwSRi0YfgF92mUiiRUqDc507O
AgNZgbITc0SPL/Gp2wVixTlOMx0YXGBZMdZXpOzhFT2JkLvRsNVrp5zG5hcK2CO03wKrUZ9MNw4h
WAhAjt9n6FhUEZvjVk9AobCkWnyE3COovnUzn4jlfJicrLvK8PLG3oIkYBwL398FvmL9yIRi/xa2
DOcJ1OlGilz7JHrGSFxwc+MKzdRa4shEEkCferDRDrDEco4MYl9xjN+QgxJ1TWZxgid+SfbClaGe
EO+0LuV0+HOvfCUMhYOYPRZFqiereOIZSqfoY1hXVapTbm+LYqon5UjtLSKflX2QtibqfGxz3lnW
+FEztWaRWIChGm15V6ULrnKAeaTtH8CNl+l1zt3311xJrZGm7I3hAiT/vAwg4x4pfty5Bx4arZi+
QrAni9fO7JcwL7dfW0v1Dw87L76qXZXQvFIoOuVZbdYpAt4/r05y3251Xr9/1gtglyXNR3ENQ/q7
0+bzCwQo3utdMi/5H8qcjhvdLizTaQ87Kcg+ugy5XmNFWdQj7JQJN+VwzztJ7eJHyDtB6l8chA0m
CvB9UDkYZvu0OxZpmvpBNtUjrkM2+5CRyr6BsgbYJ2uvXeLrxGAjLpiSUEHRUgp9crOPmAUUzesb
OlIrza3lORKX2AOepxWI9/YPQi/1NM/EWgTUrzqNK9pl4RN2jEr1tb303TGtGRlFjnbSuwqMOMAb
qmfYHHORBgGz4SdxjYb08m3QvWvFZ+hz/pW01QZV+Be7BDHarV1ORZE9n6lu6sO28SauCIDIXAtC
guzVP3y5sixle5StiTpZr2N+NIqyocTnyJBfxvPpHZILpjkdwXgkuAyHycINv4q+O4wKofeH+MTR
Ss8eZ8OLnqJlFOPCKNP5VYTqNgZFwVA7FmJJKn29deWTncjVccHNQictoP0yCZsAyiFFPnFAnJyr
eLwT0QF3i2kcLGr6KpRmR1Yx+SouPwG5RCq+v2vR54P01+M9lpHV6NuyxDtER2cLA35VUYdyqJMv
wJsw3P3JahhoWWX0IWEvBI5padz/c9a0JZP4d0w27maaZy4WZCOU0O+yD7Ea8yGDksTzBV7Y/GfR
bBviWz053M/2c7fO+t2yFZjsbVdhXmGipjrQvjptZBzXvUqM9FyjKsHArw0F1+bbwIqIbp49UhWH
4k/gJK3wqKLhc/9Yt5DxM5zlilCLJsh1JZYy9YvRUHKmCbgv2S4EDvcUpfOzVTZEQuQbBnTet5B+
Qehzwo7L3BdmsWPmORWiOJOY0YnVU08A4fkImLYV+z/iK5HozqlHez/3U4ThvNI4XcAOJrJceGWp
zG3D7llx04W6uV80xcFsXy+IArqdMxXUb6I+v1fjPM8U13htoZS+tufi2qhysN5FdhZVNK+kjino
oQPZHsMQ8j2L21bJa6xdj54vVs1mXiOMEdPb0zvyYorz2iAsrFvx82NxZOc+A32VVwVlFpIvP96j
TOqaB9yqYmIiZU4Dz+5fpcVlltpsIPvNzydp8jWILivYzByLhu17WXAI0yNV21poo0+vrHdnqued
tGjUTKu5Ov+gBHD9D6smkcfsEUvl7ksne0kibgkar46sXlf5jjqtI5zayGmqumq+wD+BFKpzhJ+B
ztZALUNUNqFP5L4b/QSwzrbW9ntVQgfhzfW79JpZGkRZP7aMLDXg1bXjUsVen4CyBzI0dQDVT7sF
Jso5VIwYRNoRkDSekoZf9n7eprmOg1//1T4DQIgdgBL5ScwzZ7JzbwpWoQjR1/IUj7OAIw2Z/OQJ
cwUFynyYM5FEpNLUmmsQ7MDrgIHvWY/lV2UTn097C+7qLgOfnRbfcKiMvgZL/hlW0RBoMDj41o0i
Q9kgtFtXD3xHP3Sm1xj08L0+tXQYIBCbAw6MEcu9FDlJb6GGybqkcVuSmjtCkM/HZPoNCztl1gxe
AdYTZ6/g7AqUQBjqhJbeOjwUTZG0l0VLgCPRO3iZMipGs7eHPidEx+4ABl7cL++2foghVBEBYPF8
XpZ67Z4ej5NscUQ9cT/UapI0v/dzTDihu6EilELZJR12CETSnzh1ZHeRBuN6d3VKNKGOqMW6ZOa6
7YwxX45t/xnIRLqDW622o3Z9VNpF4uMcHss2cDMY41aie8Cc9iLc+kejpbPBCyzalJx/rB5pTv8y
ssuRGJW5D17Zye52fjB8sGBcsG+Hm98x8c+CwSNd/vtHTq6b6QYpGfpV1oABnFC/qRcJ9iVlX/9A
Fw4imv8ihbHd02qsckpxUMobvYNSMQMhHeC4a5A0Vp0WANzktUbv6fYx4W8Nrz8VwMVXFKDsFqC4
ARrQHtwh/cvRYagTJ0Ohhvf40aRzXrprmU6Is4T6F7L3oMGYZaXbuhvb7rOSOE1Z2NUS2W5tenBc
jQIJtERVQ/w0NdwBXaDJFHmpZflDNAZib45AAgR8cTH+MN9fElmE9wt8Da+f6dhqG0Ds64+3vXxc
0BdtTQ8VyxMgrL9G0RN4Pj80tivHEvhI9G3oOu0aMwAiJcnPugg/wv0UmrQXxmRnFNLLCox7ou7w
eEzmnMk9mTHE5V8yesR325u+A8TssUyypHD1IZq9brNRjAOD8ahs4usiOK7gmzBhSzPeDYSTbaxy
bmo0YcMhpumNjlPOzgGaV0zJQ6c4gV65QMbXF7gi/3Dz8f89yaDsjzlK29s+lIVHWoZF5w8lGaOH
ewvgY51p57MVHc6GIJwRp3KhUqE1GWsnXB+5IuHCl/60TgKwPsBAxrQuWstg0xprIrgN58u8S8XR
V7YS90rdg9eDP0KN+tVYveWYYd6mzuvzfSJ0Qe6MNOXoFzK0ceidErF+XYsKrhl6XrzyT9qTfTYU
TTqQJq6bDspcWffInz3mEfuOeBPiNV2WhqL62aTBSbTxKdfygLde3M4xoVrnIcfBocpA0VXqPhQU
JCvfYYEjR0ocao1090/dCtCqMsK1u+dYGtryQEmzX2mfaL9bQq9iA+iv1CSYCY6tDFtYQ0TE7CbE
InUXW/iGobn9mChBKK5qEJ7DovBkc3IaB06mJOubJyA1e9xM5ozvMdTLoBBlvtmS3JPQq89yhTmn
HhMPFWsMmmrp4JZ24x9+30lpZujlaDWvEVcmd4YFfWdlxFW7tG08lM35ind2AS2HZgICBhNmExLb
mTXdkMI0uv1C1KmBdpuRk5oWXWxZfXoqQepM7b9yG/jDHu5gpi6ZnvzLhDrr9PxAoDtGr1a49HGw
zMaRhd9a31Kblsa2NUN3IHDicg1m/MMBaN0Kmu5qSZ1NYl50X39V7MpimZ/TaWcf217T3wJAQdL7
bLSnizoGr4eH9c7ql21pAFUl14CQerQq1lrb40BhODUXlGz6mbLGVt+8ZirKg3WmNJsX45mM44DG
sjrlsYahSFuxAiUYHGbdMPHf0EZT0djneDLGVhM9juKfn8NTIvFEpWTxvLkb5HjWBR7MLad49ytG
ZopqPcX8dP1bePPMks83QnMavuB7Bw8DOgILhBKNZ0PpUJ+V4hNk0PS8LqwXnnk9QZvIF0vaWLEc
YR3sWPYq0R83fCH5Cvj4U6EmTzI1jiSqnHx/CAPhKPylJrAumbnQ12+cr3OLLmPKBwgGysMVgVO9
YjBUKmtT69JBYp5CaT27lTYIMNqQWi+NxC/HLqdYJj7lG8rvGgX0PuL2ctc1cLYWikmTXSgjPB5e
Zzhveyymp9QETEWUSVwjiMmXXHdEMX2D0N1t+yn8OZ5Y2K3oyyj0la6DpmRpQnSYy5VO1QZXJzuj
wcYaB+U9+iqdHlGp3fvbKy2NxGVmy+OEhFRoh/bstx2dppahZ5+UXx1qv/UKKrVIHcN3DL/iogmX
1Xw/vMQ4geDeruUcrFgfwlDTv1J2xeVQPLHgIS0Z2tmrCHE+znPCe80P4HwXvX47DCV4qHygvz2v
x+a/1xbtgLtoA9dOO6/QrSk4jtQfQOsSSLR/N3spPUxCMu1AIVWK+xrxaSSMGdvyZDzjjgwrtD4w
GJIVV8yUEgazgWOt8nOymZ9fcuhIPyCV02+xfcd5aF+lz00oGuRab0ZVg1wCeZDQULdxyzLEQPVu
TWwx4tcg+k2+Q6mSBEhC6xLOKZag2hjOWkFIoQA7MmQICVvQGAlodF4h/lPrPe0g+LP0r5V6vvo8
5An/vDIGRCOQ1dovNTF0VBOtKdqx0ifjRHgkICehsUnj3XsiRg45bt4V2+DNUKvnhkONTj6rKg9l
3vXNuOL55DjkvzB6gT8HE+KmDP7MJGysS8D8E07do3bgOvZmw8oZZ5EeSmp7lVzSTIUtInB8qpQ+
JV855AmNUmTBX+c1pu9CLISBvIC8NA26TWtB4vYvyYDM4VZe6clk1RzHevdfHxNJoAkp3I91yoJo
ooiqTuq/ONPzMO3C7grZn5tpW3iAMo/PrFMkfFbJe/aoiygazd7HrYFUf1/XlUf0Lu02eDSjYU8b
BU1U7huAk5HeliSbvdI32dAC6FtozrsH9mtCeUBMwQzy8tN170tywSjMKYYjp0xgjfoAwcdFWYM1
bVhtAZm7rcxz101H9oeyG4brkzsxrYfBx4xiQuuJ+VieVyxb7izh/RdDfpB2UFi3tNGvcpy/dln1
JCnd3l7Aw/c4Hwt+8ePoCY6ncf0fU4jswR1S//GxhVwA8D5UkoCZNVHyEH5W+nA+MoCfkP/UJZfz
cVy13QOLjXJD3r0gN1P0s7+rD1pK62O/O51GHgAIOPJpFBLXKt/P/ZBuYCbb+p/tn3/dkGYN4cn2
9Ev/cKfFUEUbzbOIzFNoH1vzL45fPv4itY2S8rrvpXhUmRV6okvwFMpxZwhILek2JJ8KdhtQph9f
lvr3TCGqjTtEjQONke6n/fYXoh70LGXixZkDHCYboEfVR6ga3z8rjudMQ4S8vdxwpYcSkQOwXQys
X7PB/eWUkZJwlb8j3GSIFHX0QvYovewzav/no03rb58/LIteZKKnnDZ3gaK9+5vPkiLKDTbTIvbn
JFf/ApbqxX5Cqcn5AyjBpK3vth2FPa/oXLIUhdWUvWzDfy66KkFYJ57NjQGxGjtN8SO2vBPBCKdY
WQpij79p+01ZVjxTJd0tiu2CMA4/s7iR7HgRv8cDA03LYLgS7ecCCcPu1iWSDsnY2tMU7x6UoAU7
OTQGPAni0fOEMMQtFJ9pdBO+BDb7FAa4bf6Vgt7Bm4irjOgOUMxEuUZYDiKPSEt26LCREdoTimTA
6PrX4SNQ4MR60D+IPB5A8AdNJkEmTZ/5H0XwSdCkTbtaGlkP/ML9+vn19QCubwlB2BS3nwpFvIPI
GG7UMuvFSHocFxlmdMXBWRpQ+H4Z3EwWvZ7y2zFlN1KE+X5tuY4eHDrTFO7eWjHrqh39GrU4PUz3
2iP2X2jPiO/1WlVhJu5DqZtpuwwZnT7LRugGYoE9WuIPEbb24IFp390edhMB+B0LKy7B8GyiZ1sl
S8Hg8hDggqzEKp9H2xMT+YVm9K20XMSj2+IMK5gVT+EfZya/ZfKuLpQWFuOh2sFRDF/RscoPfyhR
uzmGlDoKSbadpyJoM6jDCwfFy4PSpKiSw6uop5wEsi73oagaP8TsQiOY4cAijzlSeFFAAI9Bbdo5
Bpn6cCdoZFSe19LXmnEGCqb3aQbIQaZUZS4DybNpT75GXRA/An+2W4DHGD/slSxnwJWPQ8Wpbwk5
9BG0scilaa9QJPF+OPek5tEw1UWyP6aLZiV7lLw4qedFEkquGMLb3Da4UhgWBB8IhosEw+LAlCCv
xFhxvBYo/WIT6zKaFpwGs27F/Tyn5vQMSwJZYg98ojmbrWg0+iIxFT7GedYXDt9qjTe/MgQ/NY+z
1pM8fF5ytqas7F++KpKH+EaQzfQoT2hvTzs1SmixaGPVWdbA3F8XvBNNncuh/rjHLpCJsQS8cGhR
bXo02WQ3mxdX+75s2ZJ26wV/P3qclG5vL5ZFkUoQwV/Vo5spGfof6RgzhD7xtTkPOfs/W9FNk5gj
lUCHpQ/Y8WNYqbVk3HYhNkQphHuYOEdWQG7yJwt/t4fu+G2I/cvRwZNatEX7GdSeG1GiOmFxQDcj
8z4Sg0xeu1Q9o9eW9oLnLJnrXneAxUGNwUEmh+kwC0bydg/r3UUxNiHsw2L2Xmt8V589B4A/kSkg
JvPomXQJbDl5CYu+RqFBx0I5VXSdU9ODIpWOLtXqwXF1VmY9hISTQlOuoPMQOgGws4v8y57aioE8
FyST0N2Fn9Sb9cWinM6/bFsFrdtDXkEWXkyg+j6C4Hwh26GnrKuwg+5OXuDpGJCRNQUaup4j/hO3
QmMLj3BhOCqxbl1p9h5HpPkMEFv9evxEg4SaDa4T9AMgLsGgEahp6sWkRF1+C9B/sl8fUqBv/x6q
73AccUIckhFenISicCG59ltKhAo9awFYFcsAfdJ31MYlZUGCs2hhWKnYUBYNteRUSJQwzIb4RB+y
Jy443eOXhkIxBPoIeT/sEbEz1f02ByTQF8c5n/rjsLIHzK5+jgS9k1Obcl0idi5al5bXxJtB3OOg
YYbIOZ3JXdtkO3Tx1WQsJrdPyZZrWwFcbfGOOIagd1lJsAQ0Fi7o1a5zSUG/BtNHR/wN6ryXnkuf
UVE51RztHGEn8CIcB2zTHGqA2HqrCe/4+2e3vyK6WT5/YWNDS92P8YCiKntXCL7x6Mi+VfzfcQBk
lfVsxsmzgNMh7Kr82VLg/40gzMPKeMaOfbfaX099TcnDcarFdawkeRbuMc+2KStkCr/+VJlbYAW/
dQeuAVfp/cPtMFBXWrz1U6KE5LStc3gZV+YLxGxHyiB2qWNn5mSl8dqp/c9RUcIcKHha+iZ6u7Qm
VDWG6LNjrlVl8snY5WkkoWJirjNzgzUQRMS+FWjBQ10gyaoJSUoQxHGexJNODqVSzKGioTAaID8K
xW8eP1M11dnoj6BU4kR88oQlJ0H/6x9XtnJC/s/ZGmzlDUq1H+1gpodywK1DoevH19VVGcOVT6nz
ttn6poFO+hajXqyguDheNb9NwrDimKtF2ZcqNk8r1uZZqOemPBUUHlQ/sExi2Z6UWOmXseGRjy4J
B/AjOj5+KvzXgREOGdDgd4C3L2lXQZeV6Jm0ZDA1YIL4DKw1Q+dcDgoleiB39hhCLaFIY2eAp+jt
iBh9CHSJydnZ5ct0s8NblUqp9U92C215jh38fcFDnZcRpJ32rPcflOZUMuoxvbYy02haCJTlR3YV
iHZ/k+uf2cBSYPMPnop9nT/kRnbmGiAAMuzMuRb3Vb27vcVzF3zGVx4Xjk2RPzaBAD+mbJMOBCId
Cy6i9GMQQrDAMmdO76/xgRkrCwLh2EY0Tip8dxe5/jaQx5nIRAQk8FvCZdvuXbwgfKG4AKoAU+is
fOJ9S4j0X3Tix0rlDfOXkSMLkrPzg+IQ4GSdQFDp5RZtOyjc2vRUgl2i5zQhmHwiyEawBg96XuZK
/k+RtIj5fswZ24wBsZmyB+RnHFKaeR2Otxpjn3WER2Hg3NkFm47BlyhV9ZuB1tC6KCvl7X2Y71b/
MSiAP4KMpgaQXStZ+2KHM3awCR4gzpGod0pPnXaOm4LcG7r1zl6qgdtKm55cLis4u88oCwv2+lwC
o6rUg9m9/RxcOGNVrkVBdi2y+A5gg5K58PMOy3rtgvtHIGDMa5+jgK8EXjxwx/C+1ujVsyJA7UF4
oCChRauM4TY8R5GI3GzMKNoYrMGMc1P29QRxWzS4c5tgHoJoWFX5vsArglO+hsFUqbQOvudZfMs4
yDZ+LAgXLJMhNBKXaDegQV8trjfKISbLeg5WoaWBoGaABZoHA0DY9MCTfXblvYoqUU6aQUTVAtAN
avAEw1iLQ1Iw1YN2wMene8hl/9L7LZs/2VTcXT3Ss/O7FaSYt1Zlgc2hfTF9Z5l5VtfFT0o03mwG
cXScXq0jgZlG17tEShTXYX6AnQiJHa1GFr2SGUh/TfWwj4Tmwx9qmWFRWsDvCgqeycm/rdC7Q8zq
WvM/9CwHLMfpDpFct5LXtSppzOXlKt54W27guIx8tjimFHn97b/Ht4BZLiPPNwKq8OTrN91c8swE
vzCHHLQfd6h7F+rjxtg79NAvcTPCXpHkHtOeD/B01rbCWLsol5gdUrnYdvoZ9dXqQJK0yy2d3r8/
It3/qQ+ZA55cjKile9NhV/kDs9M2/tZClRgYsa9L5jWnWkxOvGvC97BtN4BJXPZkPqUPq3jPkluD
PLMwngPzDkP9uFIcUiSICUPkwEycbuMDY+3AwBBr8lN/yPZemYsSeE50Z6FHyLE7Aph5u3OQv1mv
sx2i63OLxASFe0jemixfNUb6N/RNsJMqQIpx/Ti+NRvTnKOWy0siUyOEdClxzWPoSlJvqojjoEVO
gIfVwbJ0Obj9xM6BfJi4FUdagtSMEy5u3DG3le4xEE2H2hK9qB1DIuzrMNhBuZtsphzZOckrkUrQ
0cEtWK9Sf1Ve8WOuQUvs37zhBn8SQBrTiK1PMBdoesmCMl8kOmHuFBlO/uISF/jR9dU3uo9s17TA
zGNeAfQISzPSgOeZeiLVzaTAt7e+ciQkC4oopxJgpgaF9mNvvNXwCXgDSqhd1xbW9oer5fKnD95r
LoDU891gXeAm+4BvgsoIeDOAmDXYD9/yqg8ue2Z5kGVSxd9zvgWUCXIB78GAt+g1E93WPZ+Lz/IK
ofnZT6JYYzNk9Zu2SNvQ/efuDxHAdsNH8q6Cy9IPnrewmLD9HcaWhmH2LNNm7Bp5dT48gVnTkCf7
h2sTxH82F9g5ZomVlL78rUAJ1znrJgsmEsGde4zhwzNo+2E44DKfVydaVJihsJtkgZ6Va88WPmf/
ZiEYYGMIZoCvxoe90TsbRfv8VaRdeFkBxsTamqOiGOf7dIGtL2BimgMsoET6uuLA1spLqkVNWGft
sqzrABop4UC0LofI0zrslzzr34fPMYuY/qt8MPzu7xyj94HxnzX/0Mvr53IGWLN91rK2UGiRVU2B
oKhXkF3XfsvzLwpYZMGugIorp4rIh1s9mD04IEodhtMEYRp4ghYWcDtsYVpZsYbIsraaEFDaOG9N
vVLa7G/AAABkDr9oSY0PC8AIQL/JOKPEIISyd7ACdpaidyKeKkVdnqrSlgHeb5so9cT4jdciVpwK
aPFTi/Hy4gq7dDoHbK547hV8rL4pogWJfSZAf+1H4g7gF0KNeFC31tC9FuSDGTJsErATyDL13pwm
VAcZFFCEpCC8oCQr0P+irzcZuxRqR7Oxtt5YkkIuvpsPs+71rdffZzzxmuwNJcqTwJtf95fLxC6P
V6wTLutqRk3cEVP8xwzLQXtD0nMLjQGe2lxFXhKeccVXRAuKXpYf6sqcPvG+k5wVhkMmwfYY5IdX
ZKGiTJ7z+sOiGyCBCplfT40bzpop7WIi3f2FNRfl9MQb7KtdCw0sYm8cVzqYzGb2OMqnoChaUsGv
bARjJYOlNiBocqLqOoPLmfyMXFtcWHa70PnMlnTGlKiQMk7mWRKXlfb3E+cGELeFc58VfKPff3fL
v/hJoXJ9kWYKoTfo7XqBhhE1WEiAWP8ut11Wn9yEqPxEr3351BfmCDMjdfBUqCRt3UAyASFEXbYj
v7wV9H46rGeXBhjz0DxLQst1r4sYxjzIJCCOVGorKcg7IEbRqWdy6i3oqhhF3/g09mwkcE4nQOaK
m7gwQ8OBhVIGKFrBTLtLAkVPmp6slSsdiHr/16ByRYUUbTFudSdNogoNMiccKFAbgSOAp65KkyPD
VbqyXwdhJFw6b22a2FgrJMKq8ZzGYJ1zvI/CpzDT1KNc61ZI4J59zXVy6xRm1zctxbIsC7qM02zE
NFXFFsTDXmx1q8b97OZjk31ZSFuPp/gYgV8MY3/Mcbzpl0w91+UlP1ix30Y4Ql0hxNm0csESrC5a
2EQqtl+LW3fBa6pCHivmZwOcn51wK0IA+XxS7v8RYlkPXNeXwyWrNb2OtUYQNguUOJxhY5r3WgY8
PHNMrfqyHkGQSkyVa72WGBvrqB2800Vjrzrf1V17aqjTFaAYVxOeV1tXOdsys7U6E7qvi1XNuJrI
9PfhK2Bp1qlaZgWjO+9mt6oNfPgqevXIUQvTwrzbkqsDIFndO43sUY0uhVhL9j13LCvCq2pdQ8uN
KnQzai5vyvZCGULOerZ9ZFGpv6ROixWk5kbEFnrsudGoxtPyr5s39bSM+EkWiqi1EdC+1XwUJeoI
IfDlJuRgNmlx54KotDitNJVjszVM9TVGoCIyhZVehSBxmsGQfV2R+rQXqVn7+h5erpZMIpgagG+7
d9jpjtraggpnIffwG/xE0TMF+0mFtP5giLD7HD0sxfBwLZVBSuSlKUDwnYQVgf0eKL2KTqNFeJKW
A/qIke6WHuJLm77D8wgVj8dnKzsubY+gjYsjTjFanhuohVG80gDLTyaaH3wBuYnF9gFz/1od40Gp
2AZ+3YLJdzgiMj5oTIDOXqfF22U7rHd9QU9izcppXc0Jtwe4znS1GGZ31KYSWIAwo/3pqgEqguNk
2GgT4ckP1RtZ8+Bx6oG1evJ6CUDoRqhSfOorm82UGv+clGsqyKR2RgAeB09e0+S3w2FKSNz9UNIu
IlV95lV2i4MhUbZ8RLVGW60WrvyeOiv9eVL29YplvNLZ+5vUAitHRX98w+8O6aDW5bna7HgesGyn
7RGwA13LnrbzGTILH9ziaavuV3dYrF62f8YsDgBRlpniPPbOQ4L6QjwBiZe5T47ZfaUnaoimpPGP
jvvhxq0q+lyp9kpWKtiIruSetztk8ofBGHTFgit8sh8efyM19fdvN9wAabl8uVvmTRtduAnE+Lfj
8H+rUe88Ntod0guJpDJdUXkc01YetMNaULfrcpCcXtDLesea6tuhnl3T5hqJAo06sJVCm87fEvl6
T0iyn0bnUvkFWKCZM62NeQ7TtdZVuoQUNc80GR6cbQ+GV7faNbhK19Qi3D7uJFu/Ow6zI/jlX5WC
59GCMEdfRpkii3Va3pUrj/FrpQc2RkhleGaIxEHNvhhxJR5KBtJJB7zu8pcyu1Cwv/17Rfi0x+wa
/o0KywR0oUIbL6hyr5+Vlm+/qvWmwBKjJaFD88K5mNBgQiiZcNpTlC2lccgUcQK25rLj3qWREJ+g
9IEMnGmu2LisvW9RvTJwsSjjg7HN53tyZM31PES/S8bcN/9dFwWR3byAJkZofssB3ULqkndZ17Yf
Y1AYEpzbmTJ4mleJPdUt0hyvAhq0v1V5qE3di081DbW37SA7OpY1w7l++8d+RDSY85zZd1K6Pcv7
/iXcrYJ042/sxy13bGIVJu5rC927fW2K7BNCa27Lnl9o3/kEvWGN+JHQAcU27o2jIlg+cO0R9p2q
vLNRVEOD1AJLnr5ddsR0i41cDtbZxTl2E4IFvZcFB+/qzGvSgxJkzWWIPe1LQK+wRMqaNPA1x//w
4fBei37+ixwFM9+pKZlu0GwMVWIicaCSkqqLPE1tyDWJT0j2tAHqu+dQ4tesSB8BQ7Ytz+CTuZTg
goyAVYHZ7VXDR1peqXybEZ8dW7D8eUfOBzaZoWmRMSFNdoMvvpXi8w2kwtr6RCUcLveiYD7iF2oL
rSjXxSZy15nRJ+F/LEYHRy80svQkB3gTYvz6zEwrxeqdhMQSo9Gq+FDMY3Zn8w7yehffhXqbpvvf
tZMjV3BNWxzhrhbsqQCzFoipkaGvYEePeeEGJxA4D2pKpGNS4/rDAiT9g/A06oqhG97e0isQ74Jt
YpP+QLpYPTZzUaSXI0QHVpfNX6bCAj1kyy9o/Sw8v4LK79Bp4o6UvlpE4ZwarrKHu5kUtkK4guWh
fUmZiWnkBhIXLaI+z6NpGdBriseCBJG/I3Fbo+ASN+ueh0Blf7OEO3AohCazRQzOHTUmm8SUBWYm
UBGv7Rax+hnX+3EnLXTZyuzvvuagoeqX0z+hSo5vWywriKTnD62Z/PwzzTOshcKyHQSXGc9vjVyj
CNeRZlfYyplHrrHHpK6n5Aifc0HzXFhpJXHHuiqj1GamDL/ljNrsNuGfIayBNsoZ/DQ56w0qDxtW
UEJrUH58qvJR2A4uEV66q9IVPnpv7Po+bHOM7eGMCzuDG/K4CmgBBMhLMkauCDF5HanabDsz5Gmp
zszEPeUiXqGRIqXVvCFG6J+hyNHfZhhFz6hhRYnd9oRNv0dUXV8cBbjDDLUIFGoR+yrLG2/3TL/u
bSP1MsDialfZ7HmqttkPKR8j8SzY8thGnB0edbLctyEKOPG1Nl+mHRyNtbmPOSS5qp08t44Gamor
tFqyWTT24ZTz0RzNE2aXgfcxGda28rDa+9JTJcwAejiUN55HPkF10fEjdadSLxZxu9tFZhfXh2AR
MKYsLwOA6eDNKVpOUdIe65IhUm+1T5HEGK1c6tDbkyY0RW1uLJlzr9FoYLZBgMCcdkRkHveF5Rig
yBnVbjeAlTRgyNYoPcmfFw7FF7oFZVEtGFc7dXT5/kDuVJ/ubfFL+Af+mTTtv/0c7ARfTdRqubSN
kKuxjZ1vK5jyGZmIckiiRlxPCre4FRnOnL3BOiCnu2ijXyHG+9oy83EibCcyXN2Pjyhyo2De6GcZ
RclImO+CY+42xU4Bq85+0XJOP0YrdnjjxYN9BlJphld5E5DEaU/e8tLo4v9H9rdAUb4JN1AoSVfB
/UXkpkAWgXUFQkA3/6zZxQ9bxXPGkRAXE8/5VphzZtrExVDy9QcwewgnRDErr9blbm7B26Rz2Tke
6CC/6V4EEXEO9VtM2vvC7p99vNs2OmMibEXnBOfcLlWl9SmwDw38315fhUiEyejQ8mMwUnRfPHBL
Vmx8knBGdQFzx5A93TL0MGPj40U5aGbqkILbuHSk7hiSp10nXfEJxfQPnnjvExspfrh3oTjO7CNM
wJey6/MojzYByCwxoHRgFi+IAcZb9AyKKvS3mPP77A8pxKknG7kM55qHZ66Qh0uhuU4MuoWOn3S1
+KA5xIYavPs27tU+FxhRcbo+4N8CVymT7LggCC/EKepp03irMVwUqCMwvo3g2tRmArMRkT2aIm+O
ro/txpG2tVxtfp2GZx2d2rJ7XbUj55O6PyxrjRDeNFLLoBKRZTGvZwNanVEW632UrnwfPJAZcEFw
hx7CSoPyd22+oquGjgSH8T+oLiBZqoFPlrsV9DKwRn+Fbt/Dn7Cti6sMaL7USNqOFc58hQVsRWeT
ZBW4KkzWJQH0drid2815wS4EZN+/JSTTrRY4+vo4dWpqYORXyAIsW1qt8yO0d22hX+oT4ClVW7Zm
PX4YprDtrwpw5hy6Oc14zz9WyxYbE/hd9S87A9efnO1Mxl+v2XN/vDqUMXkovXWN21L6BnSAJbPL
dg0ArlYUA+z4kRWIpMl5k1g8iqrPURY7JgY+kQfwrcWUYRblz2xwq1LulKo42FVoi7vopJNrmfBM
RIgHmGZ9LrqxasQqBovJv6jUcHgL31MSfQfwh9QsQlpQIvrU/X0V1/Va6ABdRFOLmhH5prqLYJWJ
XPwMFVbRm725VzvQh8wc7My4UfUWheuoutftYmMQ01XrKdwVBzHOMhEDbPOHB3zyEs9lX62/SBrI
MFj4mWCXi/BDInIIlxoGEc1YiXkQA2LvitkmRxcKtLPK2q8UPTu4d6s0KVD3/xKsLRTnoO8ohVmf
g6cV6iKJtC3tA2OiN6RwiEhu0z2uo7ApDPgpKuniq8rzpW128J6Z8PWDjEisOTi2RpofiIGlxbf8
doY7YD4QSL8DXMcpg4xmZj3JYcX2Ck+00PJkVXUcMDXGRZtJVbt84tt5pEXMpwr7Zw22M7+c2y2y
syQYTt8wFqqoOXEx76USCEFpKuKnYvu12hqKfAfPNWpMU421BQS4K2ESl2uORfj7IG15hV+FOt7C
s7MHTIM/PIwxwQa/oYA43Dd/177qHLmzkkt8DxRS0M/qK78gLI+z+LVeswkOkUZPKQCSdLV6jHcE
aewY5nzFil/mcu2TrLT3UxIFlhCP5ZGtK2djXINnF135q93m2j43Q7ZoOUfVvS43sa0F6QMVrpEq
L7ibHoQf6eNiqTBYTqcrHRwFdQPT7UDE9pDhLawoeve2iCNi7+5/nY2VSCgUaxzN+S2BC2emZFX0
a1FTcRv6CPdgGKgAA+0l38sE0O0U3r4m7UXJYxWUx3iQic5/MChbWI2iUwHByWCs8Xu2/Yb7FaD1
hSqXZKiBTJtltac7lCBXmSoj0fJ/kk4vOxJUkeEoHs9k4z6GpNY+ZpkgduVIa9g49EIkcenolONI
6v/Tr4n6VvxzBiMRJslIamb3AM4fKBSch3kGlOUd51mra5z4Mx9Zcy4EPmxXJRuczMEVTO1dZfLu
n4MFTasq2LC0wAxncrRAnDsGJb877FbFoYN5jc+Hn52UHqkMHEbTfr/dZxABEo8bl4JhxydWIk49
z6z+K3U2id4VWDfcR+AjhGlaNFKjK3XMxa7lNAHbHKzawHjDihDmU9ZohoEyK2xFf54fFsJVJ3Vz
6bHUKF0zffbM93fcfAaqxOXh3Yr5UkVnOExZHqXhNGmZHHo790qj2ZFjp8z9dxmu403AJeKBikKb
P4iWCjk8ZDhZPcfnQw3a2vnxc5VvI4eckOifhBqZ4wX9xsp+J55ObzQcWZuBNCf5HmF03/lCmv8l
J3kYULs21DIt0FMMJ2nt1DdFDHmE95rAxPwlp2OmXZrWJ8Ack0B0Dz3SLq+UoCBfX/G+JqXxBnsN
ButODxiM1eT6w4aLI+kQlRXQyZ3SFDMAFqo+05AQDXxqYRZyFPRZGVw/d6iVcRtpgBvJ25q9QHrf
8PF+YHTnXrimDew8hUjuqZa6aYo8NTFFyPOewze2GDd139qSHqrEMjoTxO7yGQ37ncfnbw28KkIF
Zqt902h3y8tGusgKo/Fk0hk63qxS1nJ1xRYKofSAUKLtPIHOCIviyDCQl648AXsCBWfPxQ3ly8+W
jCe1u/xwUoOxa42R/fY6+ddeR08xXHap1m7GgMiNPKClwyxn3det1+xFYItGeNQEDecoKWjs32sX
sVLr/v7o8Ca15QmQs8YXnZG5wi5NyDQLUASWCItLYuHJqqkZ350qBpK6oNZavZ8kfusvpCWnePrW
se2wgi5RKkc4AhBa+JIzcpjDBUoTvSF6l+3+xO4W5l21gCZvO3zBFcaMK9fHNnqDYTJkBAgmcTRa
UFHdOtPSbV54Jif7cyfGFGeilastS0d8btaQCkg57YrfDCMkpdKlbUjiTRnne1Y4RChx5iOhgfGR
yM3CYkBSa9d+QV8eZCj3KDMhllTjeFVucHeUl3masIOTcDFK4cPfC0MNO+QubnRDYlJ/0e/dHg/V
tYOXN6xTXK+bC1ux6Oyz7oskHBsFQgCy/0sT1zRmpns96a7p36OfCFQhtxRAhi6ly3GMjbJbo3Ho
qMUc3ULYYJtZoJHDWFI5GH0eqBId5TopDE1h6r9TNNpciQVXLwUYkhuvJs2cKXWAIaUfci13GHPq
MATQG7CLq5xygZk8L5gFAg/S+Y/WAJFAEMpVutFtxvJxTeqBVpev9I7/pQI8PTBPnqHqakNAFPa+
td7riytitg1e7B8Awfy98vMF3w+0iT5hB1XSpae53SSZKQ0sujtb7g3WxmjBQBmBk3WHhPhVV+Ol
PhzNQHqCvJqNA5czvH+SiK/8Ll8EMhSdUYof0OHLtzX3N9pOBumQaSTHFDiLb1gpiiiXGUNSMEst
ao/NxqGdzzFyQKLFCIb0RTXz3y/MGzln8p/11AM7vYh3cqcvFmpyrInvN6cJ0J7QEEILjA47vQY7
YV0KWMvkuEQYQzTk3RK8KhMh2utB1s+/41ag9Ruj6z0V71e1H6UwvJUl1t4SMvZ7o8UNXugYZzD1
tNtgkSF0w0e9VuIFySHfNUagdhggfqRfq99H/zg4tGv46ePhr+N7W56nyEFxp2GDWdEVMqrPPMFE
3kpRh3UoHzRMCQLhwbCc2hSuGm8mMOfDCn5zjZLd0Z88khMNSUbKGop54HnH0Oy4WZmycdcgppe8
fXAka+FLSt7H05SiLB1vSMcQpMknjLzfX1nm/CNXRUhlmc0DCJvnDUohRN1ryaEfec85+01ds18k
Yq14Ml+ZkE2U11NBlURV93goMcYKWtrwReJPHfmzQ6Z9u4RDGfvaLx65/Be+0i3FQk6lrvk0AM2o
2pivOS17zqXcN7GwujX9f7xox64oIYQv8C2GjmDd6MR2IdOO3nZ2iw0DRQ3geoFu9R7a0sRQXRtD
3yB51bCyLM7Yb8UXRfMWgbxXf39+aX88P1lxjeDBldhOrXUEYjlxDaKOgd8gI2ze3trIsePKGEUm
bzM62QYgpJGe2h2xUGwIJqKgn6PHHPkSeQB/KrbPICq2tQ7QwsRIvaZI2TGjDAJRoiwigApdjcme
6lSXPFiJiRphPUu97jjTYEP7bSiVTANYQygAaH+woOaM4TJMBQPoOv8jN0+IurWP1Tb10QFOs0D9
g3OscgWJ5NMEwW/o5KZUAlh1rfUi/v+a9g5V1OPfDsndJfOkrh70vSfP81XMy+K8T0yKQ/MYdBby
biX8eB/g8zYUyZvtQAUpq3nUhIIyT8Ne3gkfBPXLeT9N0M5YYAxjPy+BTA7oR23268JQh0iOyvfB
6BVv8KMm47fQBHuiOycf85wal1IQWYp2/nioSNmKXSXzkWdAjafllDp6DUGGaJXxKFthNX+lQFUR
UPZ96PiEds7ZVH9Zxs9e40oghdg+A+DemCIDcOji68zfEghiN+5OugJBUVzb649SKJCdhRum2cQ6
4cKFXULDBHL/AsAFSgi8HfEQJx2jNsBzM0YDrlKoiTl06KyXkSBTJEEHPIgOaE6JT284vgVtvZId
Dse/HsfeD0ByRyu0tNPfxJRq7RD3CABe5+4q8s06mUhZVZ18Ys1+FCEqjLAWWhH9O+sbE/idC9DK
novspLGHCt4+lhWBi+B+Yuhn+wcnzG16IPApN2WWdvMz98H8GqrK8l4LtEVT94rHzBTDlvzXJJHW
VSAe1usUQaFt3VWMO1mTWxLFtB9eTSJzzHIGRv3dd1a5cSlHthZ/daxcNGlJaglbFwbdi1RqCBej
YNM2uNXz1rIHaBpl37rFvI3e29ylKNwR4kwBagC/22tm7Z7NCpt3v/jXTCATiu/gRy4+5nVjV7LB
baNELfzH8GfXFRtfN34mEDg/8PejzUDGr8Rs/trCguO49aJhdAcCp5EJ03rbkAywdeUh89Jq8Y+8
bIQzyYHxX/pWhra0exbLtV8rvi7bv0syRLcwwyaGNRPvLIdHLgV2jIv0axLzIZG6gkzc/XD1ZblI
3lHHmfbeir7nZMwyJrB1ZEzYgNcEMiI5C7tvcDGdK5ckWnXfr3nl1GVWGjcx6Jy83GmYDYmGw+YN
j+MnEMuVH+Pin/igMPRY/37VBHfP5ezZLV54lEDxJwbWMQ2GwEPXFhOI/XcdGU5ykqzlVY0EORIA
OLh96Op1pwu6YKG3TFvZSZcfPksczb7jFl2lUy43Y5lsteAZIeMaFjtSXYOpLSZHHZotRx4lrld9
xh7VCI/rngRxU7ka1a+2iqSjoaqJS7wyVX8/oVJ621x1+rvobthXCyJrM2+9xD4dTONpnlzx5+aw
0Dyf0OLYu+uGi+MNVX/q5UMJmXJUcp98tqcLWhps3blP/majf7onvhMEsuOm1foLJ3T05yoEK1Wa
RTO2gXZSESqpItqjo2DDgkFnvqoZKmqwy6swZBvWPeesjGRoztLCA7/H0LDg7QVzv0qIY+ZU2TuC
hbhhHTgy3mrOvz+pyg11e98CMJZCQlIqDHht75qbu8+nTGT5KYDK+iLEseRuQvdY0qBXiPjpnHpb
NpBZ6StroSjibwXZdKxQVzjNFhktWiNF4jjEvFlR5JcIdWXy0uZBHfajt4a6pml0C80pcsjNExCS
9qEJUwXRFlpZktrr058/UfBW/ebzb/yBCGngQvWN39LExdeE2RAT4jyDBQJgN/yd5pxeGACfw90/
RBB2/R0u7sJpv4vwi2gXXQLO5hpREN4QOVeoPOwLzYjm/yRTf51jjoEdKK1vc6KSCJcfTx8SpZTt
p0L5zT8HxghBbUrrbTPz8Q9aVqWIQdjdW/H7bTnrHZRBkxaWlyIqH2SXQxr1gmM2tTHL8xYyIlkf
nWvyV9Ksj5zJRqx2EGH7iJECTwofHsVqqcBDMRtmcz8KHWb2cSeK9UrYeRZdcnYEbnfxeZ1lF0ja
Q5aJjhbIEeZPwrHFCMKJo5ezy2KTHRjkDYHSO12xf+XUqQQKRnG8c/BBhywkWpC04ipxYSjyDv2n
djkuyuSHruZKZXj1CoTW76wpVAEu36/pYcO+jiSRo7eCA9rXvofku0eZiueYzofyAn82OBLiZZad
MM8f6d+BXeExXuXTUPYnlYwndCc+LE60FHhuDpDv7b3PwSfX1U5YeYIIJZrUEIuHGn2ptO0zXTQ/
N6AbecVxfCT5/F4f93JXqKsfOYZkO9xSGQh5V0txYuFIWWA0+ZmkGnMZdH1qjXTWqV6Azf2XHeuN
aXtAxfUxoZz01QonWq8KeAfQPu6bI3vhnVhoUZTlJF0exqe8e4DT9admEtVNppMU3U11sIPWUvhf
mL1n0tZ/hwRQGD9YEl6SV36lVtoDOn6+0kIhcADJ46oKjbnpgE6w9IQtZcrbynkqUUjCDxqo4g3J
E1axwAxUw1p4uceG2jlae3q1ij7XjWqbhN4m/iJ7iIBD8o6EKS+7E5HoLPs6mwTBYNldlmJoWiTR
N6u7wqU0xWl0SIDqja9vazxpSvcdk0S9YuL/23TtSbKXHgfDgtkdf5H7qcmgMclKVUvIDDaBcuSK
43Uhb2kwRuaSTGpcd/O14/yCIyQ+ddsGqUmCdVuENnW7c+GQwke/zyiaxC+7i1r5i/o69W/HMX4R
fUV9yscWV7ufZljhOq66OKL4OUieJQK3veJ76R3z1D8Dus4aVAs+NfJpK8MrTmEPzZa0r2q3rs6t
2m0kBfdeYkYNYMrPZ9qaw975rdqxCOLOx1hBtcjOjIRVAOp5Ur8/YEmUOyQGEHl0aRNpxvEcGJke
tthf+t1lXwYK3cyebNsL7JyIYajWO81VYBy5CJOKkm2YdvJ1fu8U/UViiY7t00kmii9CSbWxfyjP
m2D1K8N4D4C4iucOrSAaetyjXsS06R4XXSVnZHfwNIwfxeVZCRlvaFe1XEPdSke9d6hWrO2XVGIa
jjR3uzSrEOwBGUBZcXkDXPEUNyiZIOk1TeFSBHQXAE7ryV99vtjKTzo4gRswnCA3ZH9Bogj9Bxnn
lkh35zLkY4+cwjeEvvW1Qk2Cz+zZ3JVM0WUDCXSFXMBCniK50Qs1jmeo0Y3j3HdTHBC1JxKvKCWx
dwIZ2UZLJFqhIY+TTcjkZZottHhuPjO/kRiEyNZD8kruNg4V4nZ8IR3HAOOqiVeNgYl2E6wkFd6Q
4at/uaun4cwQyKzdlMAu2AI32pCN8+s/7ADlVCQEdVCu8kS4UlyDFHJP+2ZlVc1uME+b9wJMc8H/
Mq/4vxglu6vxQvxM5saxfRLaPwdbDYQsCP2WgfMmTzfrg/q94n2B/wS1xYFGyYL2kx7PStJ0YtlA
zbKIFauWnmMzXdDFWfnH3PjjUKaPVCzaa7iD7AsXtMFag0tqUbICsfs5mByibkL4N4vYI4+1glYG
C0+wA1YgamFOmYOR/inDk18XzeNTNbsnMBgOeZ5jWMNScZ3Si8u+Ydx62iJKpTdpRN8b27iAQD9X
MsgHoZEuZR1yqilKNUToAY1wmGY/7u3KKi9CIGGFJ2YJgRrLA8Xex8BDL4sMKu5sKkTyz01TCqMh
ziyhPEdKDkrAC+vEtowM1QJaU1voz2uhvS8PJj91MhW2DdMY0BY6hq9vlfJVpghS3LmniOGd4TC/
zrLsVuIjjqQ/4ag7poqPxwcOzk1olUP9sJTtJ6woYr+R4PheWS+UUSD6cjbh/By4aMJnCpsTB2Xx
0clo89ZD4zgZUErxbBUmACtFxgEZM3sk7CUjyWk8Am7R6AJ4hT/BDfM1ya0Nt5oKQo0d/0dFaq60
akGL4r1nPiCZeYkDhhjxlSVSOC6jcba8jCqG3yJMnPzUZ9RwD6GCnbsafnK/2o3jFdwiL0E0TR8h
I9wrH1iKrKKJME5l7iFglIXqbTP7dv/82MgyxeKGrWokdNgphInW1QNIHAdJuTkVcDS1Do3pHmZl
UouNt5eh53JYXL3uvyl2Uf1YiK7g62cxeB34r4LNvqaxldMC95OhRVoNDZX2u3kC69o9mEuTqF0Z
bmBO7/50F/KrTWoSxABmgcmb9XHBKx3UHQ9ia5Nh1J6LHSJL/Y1bwk37q03Bp11cxD8P4f3rTVsM
WStyi96F4HWbIj0v0lgkrWMaowyFQu8qGcb52rBuzoQoYUHgLKjADGs8xiaKdOKCWCG/D9+SiKpx
ZlQwLaoll+LsbyNXKtrjOGzbl8w+IEi8wQ2V0Kz67PUPlt4ckvRjmFb4Lqw0+lIHigSF67PCFWAM
V/k0+xemwjOVGsBgEUCSLiRg6u+Pn6ry+Ckv5QJ6bvkPC2l7IG7i/4cORyfeZLV5/frSAt5pPCUc
vMgyOYKzbKpNbzR65wgvXjkIFYXA7yZRVPVM10swOepxXqxQdiiUyUmxyH6g21k1luftUjfgA1Dt
osGc/Ni0YRGFYcghUCkhco4ucdai2g0QQ9l6tI8LE9TZ5Z+LWB4ZTzQ8c72MUBz6NUpnnVXdr3ni
hoTr9V/NG28X96WG/e8YUxOOqIsjpSGFpPhxzUocvqAG6or0C5Vk5vfGGYZBQyy9Z6EBT82L1/jB
xxQNES3D5ykz7Gnek7ZEXH9lEpCNppODfggkhzyWEq1UjjCMDCeWFAUhz3gHTBl8HqhvudTRtQDD
clzDZsrE6e2Qc0rvq+PX7HQ69hj75SVWGVaIk7RPXs4t2eRikckkowtQ4zp8AuOpPfHlaoIdRBXe
6mkEeEZRoaFPnL+JshYhapq6Y0qxj2+YNRESpg5SH3+fuW/+BqK380VA3WsK7d2i9lOoaY6EjkgD
dwA0nvEmwPzRPdzllQAlqZLG4kOf8dx5fvO1TYFu70nOlB3zpHehQ9QsSLbIU4M8Nw7prkRuVFQH
PKsWD5zsvaT1lDPDJN+EqpFp9PuLZYC0k3A1HiXiRhAuuEp+Y3iiMJJdlNpaBkR1Pn+bVU9yyEIf
YK1f8zvwphbeim1gcjmkw0MPrF92LYH6l+jWh7EuMGfwefAqVHa8tCELQNocUYadXlqJ0uLRGoQz
HqYLd5tl5I64N4FTY2wry/L1f1ZBlunKwXpBtPR7mIeNmKsn7sRznPAUZm4ZjzrVTtC9T1LfDnJh
1W+kzjpCReKYlSMfqbzg5kstRC5VrQaWjcFdNKqWFZFM/J8lTlHUsfhKzssgNHdxTsABkqK2IrA4
PMmoQZ1jyO7GUJRWX7+1RRQTeJim3aTzZI1oOEn1iiyiEEFe7g9PvI99HuthxmXvJsWZIg8IsgQ0
MxwlAXay/ixGS6s1uYCNS+7os1XMc8FNyYR16TyvOpMKDazaqxHUfi4CNi1btwDidxRGprW8u7/0
0Fhg/P3vBPPo+/60rr+eCyLx3O+0gW86XZ2p0SXwhokEUSIznbfU4bSnpitLCZ35jEDmaJEHqJ1Y
U4+YHXukDzaxVexntVkHv9cl/DdLSuF1yz5nxRF2pDq892f9zsBnjrvEQPHrg6owWm6Vh5Ccx/9R
rLTSlL1cjprw/VGFHJwbjNZGoYcNCcqy/6ewv7411+Fj5dMHYShATjIpjgwwyrbkJeZ+Z7JoOUr/
1D6qV1OQDqZwjPcJVWL9F/kaVtWqE8e/2fXfm0KhaBxK2aDvJqdCAXD8cXvP8FanUbXyYcSDY/K4
onxHqM9qJVW5A4RKXs2uFiXPEmUv9ZsM2wk/2rJY2ejOJffybytwzZPPPj1c58VMfTtdrOROiwub
WVMHK6tu972+huNjzu/CSHUCPNNbOP56RkOW3+tI2pR508hjOnAwXsKFmvJE/Qhov9Yit6bw4OVp
TEvYRSAv4f/uuBkHZ+hnlSNl6O1C/oU/3lUV7uzV6x0URBK+X7es/xIEj+/meHxlwjZzfdeydpq2
Z+w0rYSm0KHnOxUGjKNFzESMLW8ppE8+S24wDWPBmKytSCF9iBJVsYCymsfzqrABQH5v5+8xO3UV
slm5iYPDThD99fyP+FGn1FIii60LldkQNzhscGrsSAI2p9l9ZJxqqybLyQdhxQcDddiEszkV8o8n
55jyu4VpnVlGDfRsPHI5kfGmrT3kikePQvS1vOUNfFBF43+DKGI/pAWazayyIqMdccObCj03DfHQ
2YLn41Q1g3ZoEsv1rRN3+8EZqn7z92QFZiJ4ZaeGESK+4sx+3TIxELH6HA75qe1hP+izk/1zJFyx
FAWGaTOcjZWDAGbtiCn72Z25xkYdpmTZyJXI6ZQPHFp9+0+6z6uY+sOBZNf98pYUeyGUcRrcpmYy
hDzHleGqjc67hcc8oNA4ScJy0jvHmmiswep+QBenCd34KpLuZIkgOJ4kTy1LkQExzSEC0GvUCjbH
pjnXuwYFLTxJXnG00mUpHUqNh+urht/YqCgTn8IO+Rk6lY2oaXHp4dDy38F1vDzce+uPu/chiB2y
qccujGkfLh+U1I+wwrNAp+aCW/fqoUB4CoeUE1Vp4N9dl4uH7giH28+T89vuAfw7D44ktU55QjRQ
0IGYr3ptuYlUQW/jIFCTGj8/iiOKZmBTyfLhH7QzZLv1nAjTTNU11LpkjQ1s4N1KtM4CTUomSUxE
2KkcwDh1tHLL/uuwFCCg3VF+ZsarLR9QGUxVDr/xm6vHKEm92+ySD2EM1syMxkLwHNmgUdpjjX7A
+dnwxAXQ2XFmJyUim0zjngOk8qATO9ZErdzA+Fs+BoyD4Nb2QuPHmMqx+OVZz6dKA3SoAPwQ7BH4
q+asoMWtW6nZJSCTYYjNrm30olEAmsK9b5uDZh5ck4Ty9DjcKYwF5RCiUaIFdi5r0x905POlKc1+
YkullDJovc7hdJ8ATf53IDu1OLQYIRRHkDuz78Y1OLARF2G5f8jrhhxxWYGeElB0Nu3J7I3vh2tu
uVZKVctcowTV6lUJxe8B7r2xIELj2HT5dQ7UNUYljxvmheVrZthvuPJLfRP+p2k2xyd8XrmNeTZy
IdTU9Fa6KbDrlKux8gGJYEFD0L5yLzJQHhfs10UT5yUxZGzYAU5n3m1ZiZJnU2v1FQyrJbUaX2p4
Ecs65cPXmJIBSazEknyuWhcnr+7x8xenucZDb4M6zKHQ7TXhwOda+6ReVTsTluxXd5+k9PKXfy5m
jL78bv1LQcLZc354hl26MpA/XNWqI7x0rjJ+dOO0tVmXlyCZ5cccn+TicpBG3KBDdeeA9RqdkO5v
fSFkIfBQ1KYh2N5rDfeztFrP5iJHy25YAYL5jueQ4gMe0IY1NWpW7OAFZOTMuvVaAgcmryBfDLfp
qWHZs7H1Kzl9Qzp6uxmsceMIKsxb83unzAnWgWp7YD4KCzzfQB9qVPeZVuedYEqb1fLK5tsEMyLo
6KNmSed4mDbhb8AnpIiNiTFZ6IOhOJczqy0QEXblAb/gnm0bY6CG1yDFuUQJgyQg7pwJ54Q55zKc
tKVA1TOWQjcIG0xYWoV/l8Pa9ZY0aDczBYhTLUd77aGmxaooQLeg2ZEqLUWdAsPS/6QrR4mQSzCj
wdJEFHzRJh3QqJmPGqcNlKVNBI+7E745bChdEJUvpGoqIlRmPwopbUCoT9iKPsGM9+gK4KZYIUCr
r04OKYGb6NzOU7Vlk/7QLULYGDdfnFhjlzzu22mSKQCmSjBmOrxbYyj7mCp83Vj/izuI1+RU/zfQ
xPUN6i6gMCyQslR5MsYKtl6RDPkT8DTLFJMg5LBc8HVhNhM+jqimN4/yePY2IB1rnHNGmDin/KGV
1hLZUwNY6L6rSKRIwygrjGtrC8ooP1HfJVmzq2GYklarOZ9NKSxSTZE2Vu9EkN06ZrgTi6F36QMt
LkA+Mq2AWAJT/Nu9aJQuZa1eNePXNDg6zdyupVzYTS6pkbYIN17A3IWUO28Lgag3+4OFqWJQNLL6
pI2oxUeHwXAhZ/iduKhx4tm7ES8EbtJDnsLnJdIFDA0uEB1hgMNFeGIDx7y+jyGXTxukD/Is2fIa
5JLBiBTrQ+afwahsD4LjhWOB/3NAAOLoHuTOkh8sM+vuDnp5V/ERhIObj0KuxQMeyH8bmwpXVlhk
dThhHneCjvqltIcyjJgfrTWbBYY3Qaa7e46bPHTTjeG/QaBhqFuQuafLiEeb7ZG+0FDDIcelgJyt
I5OxjetvZS0aBG4ufKS5ZzhyF9/0lktUNmkP1mtriAD83qZQhZP12hmM1F+9VTH0U1Bem2QXYjWB
C5S0HEMLoJg5mmdu30/HIQ/S1MnZR/qv4q4CfiaMhQe2fLRepTNNzOLxFX8ZVGs6mm+7IWNdl0M6
FR4Udej1a4XruG60U3eFib05V88fuSlaN2RdqBVxDDizLNQFeWYcso7Zn6lDg51tnrtnx2RfBbu2
SY9PYKjtgY7qqlTGUl5MWnf9f1czR6FcTPKII1Fi9/rZ4LMIJE1RPpOW04cvdLqqkKSGCKZ+VuaV
dKRxxZBwYD9v1v713OM2TmZr1/nb9SwNKK+yJoEOXTLJqgpLtLjwfTje9L8F4tNHkJPex5I1ystB
tka+yrdIHsc3EV18GGjmU0K28RwXq5YzGxkOC8rYb3PjZpfDJwv5qRzxxUFSS6OanLzJk+bUjbiA
2k0zkCj/WPjy8oqSPx3qhnLXvI6iY7gI4NEL1oWIkdE2t1vebM24qxzuBqFd6nLfG3+bTv4aa+uD
orOshc3u4zjGSL282Ct5xsU78m325x8Y0pFsmGLigxdUXKRphLXemcr3a/GHt2Qvo8jyzjxE9lAH
+ES3uYh2HdqBlTyWHC6hWonKDemGLBa6FQtYGgphlTlZkrYE+t+bxUWyrM9s3M9cGyuI38rroieh
YiGCLd3aBk/okhQHj25XMGYuvVL+CkNUKR0UXuTv3Gg8zozkDVLCGIfGz5gcz383m37R/becf72V
oHHwfh/9WwqSrIdXBcQkxHTGydnmMvgfOEvmpvypZfaS9RgJ5FaaeOdmPsDgRPYAUr3E4aGs/9ml
6LOQt3D+KqI2hSsnkdR1+hI47+17YeVq3ftCLNBfs8Mfh4qAZpmR1uqQohFql8QJ3VwWLR7yoICe
X8h0L9kE4Nx3Sem/QmtK5pEflwisoEpg1FIPsgbhWUMba5KTUY/dKfYKHRJbAnvSsqz8FeWgbbe8
R8WYE6WiRKXlvE9lCUudtvnftaY1W89vlAuCo//IzH1gDDrZzZRIOhRGxW24b9BSZj7aolE5VeED
1BipTxcjVp76lxq9cq0qMFiQG6izjgBfoojS9TdIB58VQOZ/D2QWHaP3CWEd1rPDFBxnoLt51YiH
fqhbWtu3movSfkTOc8/HW1qxBdCjyrUcmQqW6KMDu+TPxG6DWk3fuLoekaJh40dC8bqED7X1GTJD
WuzYaefX88jn2Ti/fqkjei1/kkTgOrwfz7fJciDmWzsrACgZVlnB/dfq4cVYRSa0PZcZvu4wsOd8
jhcza0NSVQyiWcQetgWT2isHwrS1Kqn5s59HP/GJcsmkFQh0t8c3DHrVKu+oIXKueT5kmHN7uonk
peF4yF9MYoMDXDGKUQSIH5gsSmJ46MGouti7eKveOh8zVQ/M5U9OJ5zxJdAIzeBdru7sHGPYnkOu
c9YAZuScLNrZDQQcYjDUffmZtAepAr6bhPfK2RVGmubdyNmysxlLuaxACjYA224K8IzVjiad+YML
GN8q24jEW307HxVDXqKdnlurF7tgxyxFuJq9GLqbdWsMq6iOlNgPQ+yJw4IDd1FL8BJodrvwalAu
Fp0F/pXwnw33P4tgEGMdMzJ4J8etI/rvHz+9q4qUMJdOUikZX5WyUJ9fPQTk8wEA+W62lyQSgWDw
22AICgbAj0+nqrB9dO2OwPt3OP8Cm4dh9hlIPn9Hz7eRXLZf9GdCDxzOygefOMsWPRhjGZxXXnBF
rStReUTozquzk7kLhPfHEvf2agVUY9RGKF0q3UYaZ+N8VKn/Ieez6wMpEtcM2r3DqN5CRUOdiiBt
CWWva1nlgbNsTnykSkzrtZ/fN/sV8F3asTmUHW26SOyLDRVWYBzvPDqsCersAK6m+PrEPcjQIw1t
+k+DjznZx3Ai3n5yR+ruO5soXHFbpbsVTErc7dLOmPxz2nR4UlpqbKs9q4V5mIyjMKzv6sXlntLl
U5y6pXy8yMMT/FxQTwBPOUjKjPCh1NBL/ItLDw076oBI4eujyCw1ET4TUFZhfMdHGOtW+UsS2/Jo
fCXUlnY7HTz+qzxTsYFcX9fCbY39Batx4kPu8uGIofEC2ey77aYTdzy5vjrKTLvZyObghZXQhWJe
DDpOoAJ+5tHRXmk3DUR65ZVetj3eGa5ZdMOE3hOlHTCGsSFx2lbD0OpQhBpG7d8aBFRrUvlKSzFr
sGMvzfvOEagB5oBBU3sBf0eTwwAluR1zdM/a5fM2dO0e7eeUri3bpn6R7OIu7haQHYgeqEqVBU1p
0tMMcDpaLkRXA/NNUyxDLWrtdKfGtVgLmblj/2g0T/lkhEgplyH8yhYgRDj653kI/TW0hYDnka9w
3s9HazQM/nnm/SNtgtAOh1n6aTurCzo1r3Uu9ttjigAii0k8XPjQKvZ0euXhTy7AuBZQR6lYwcJ9
aHZMfNhyiZ9hMz/k3AJwsdIdeUS2K4c8drFSgBsT9lkP37lZaRjqvq71T+OQokFlNl9dZ+4N/n0F
ATV2/f9CmlhkZ4Pp27UEiJogX1wFiLgPWfKreOWsUVdacSa/9GHOT7Urd8f7JMp8bpigQt6CHK8C
rZEiKq8c4TpIiJqbFE/ReyKRz4ZCQdKtAlPgEKiKa7MQ/m/HcwutplDF0MKYJUlgM3MGNcEjBEHY
a3tP91aUhy0FxDuOVHyikBkmmCkKGcslYHlrP+VAXZHJQ7302Ql+GEbaz835s0yxjUmFvbI91ZC+
Pzey4f59zj3BFTaU43aW4FgibErgQypq79w2kdk0ngIYVgPHoBa+WV1VG3VbAvQDYbmHDDpbr6/9
yeWM1YGJi4XXhMUci224c6YmgVIQABy9i2Hcawx8JAQHNExHgKNsNXMfeRlV0hTUzxiLcZVGyafE
ujDr2618J6vN4U5h0GoK0q7SSbhcRPP4cUbEO+tjtclO8NRPNj1XYVbXxnf0/N7IZWRTDJqrbIGy
adOEXGVncHDi7NJxd1VCUvLfzvpISSz5hl11ADonH/kxQRGPC4RXmUs8pGVlEfEek9u8zlsY50e/
cYvwbeV7yO08GQb76yV2kjx8Uh0oGavNXVTu0w8HwV+IyuPbnFYD60VhMI1T1Xh1qP6PgkOd3P7M
0nLPDUgivChDOqEuDEXp7DnnbVKmrWa74uEDei472D0XsFXKNBsYl2iQdxcTmSHze1jWSYspqkb1
17sLR2Ubzdhl6zJq1CvY3XPI4FZpande+Yhe/RvdjAkP7aYWukxYYYPY30Lso1Tis0MCoSFNnnS8
MIfteCwvAHIawY70rC7OMdW4UddUkCs3qzCAkujhD2/N0KxCGA+7t67MlPen/avdaVw56YRhaED+
QJi15v/5ElMwzv8FZOcnTB79doRYc54PF/W+7EubBc1NetSo5SPNByOgcG6wvfOBfHEgv8vTQWs0
7ntSDAx31q8I3dT5uIUbIhY3PwYqI6yeO97gBBMqCwYvUEKnJpxa9Ixqvu1cKF+9KiN3noiMWVph
CapsBIxAhvKGEzOibVWgCDE5hmyV0J8PyopmL2MRKWN2atSH/8/Q0h1d/5r1NBOTLTYUv01XutaM
XEXtzPP60qUNh48pSgOyMPTw/U6si3s1TuO9flDrcyQ0j5pyyQziT0Vo3Cy7TNBOyNZRdn2Un63j
+1Ja+XIh6bd1tlcvkIYLZ1O3/pu+M3g9S8uLKbLvd0/25iuRjJpRbwXldsqabMimxXYnbDm5hPLU
FtAD1Psz+xW2lJt8wOpaNgzBmiVEWup/Hbnf+9ZArtJo1uYTMxWmA9f1BpezrrXc+GZfchY+5CVC
NhEOt2oCgPZZNJkg1eOHrxijMQ8jjOx1aILOVTuQkJnjkZqgrtYB9RnsJGeIVNbJEluGsHQFDYdI
8vIVoQ9a/DkM5bA1Kr97hoL0vVwqYQD+CKG/wZmB80SknU/3tj6boGeVygp4kIMq/6hAfuoJEqNY
UEOvpj8botIl0QS/sCR/Qv/OJfRVi6s9kNnN4CMHyO/AmonBYenrc6k+ukOS4p94xZGaZ8V4Ddl+
/JVXm9MK75+RWE7YQ2WFc+9RQWLWMPNcklo5IHQvzSJSVn5Htw7aVrrN+XInYo+eLmUdSRpnIkTZ
pVdVTOqpGpPsInMNpMR+6vtl1ypaQnVNcWgqrimQjPOSr9/2EjbZ6bhQvPaW9Q1+53GAWYz4B5h0
cVlBHorzmNp2+wdbpOJgNLGktagcNSu2xS2hI9W3EV2ltkr0Ir7t55Dwa86MAmH5bgz2eQOl71Tu
rhDLAT5QY5yAgYT/hqXCArRbA/821k3cEAfkd2fQh3zZHNKsBCaKy/WDFusA/U1boZqETMA/iyiz
p6LvwP7mG4jY9Q34DQ37QCes9AzQgbVFcszY0LIhBck5wUUZv+VH5X1k795ntPBFIMui6MIdKveX
X+7Or00+aEnkwdlMETYVBMJVU1s5dRZoPT9qUkF9/aLArVBrfniywUyvTc9Y0ge7IoKN2OWHoJ6d
vc/KkeUbA5rRKEr+xU2vNYqnwLynCeuqU8s29ggIq+u2rM85G3dE9dz2w1QhVuV4sfwvQ9h5sw2T
BOLmGmACTxuB67eyNniSjMRcomQtM7ijajgnlhcI7OR4oZuJGQFmOvoz3qMijOGM9iteq8rVGfjP
jwTr14GXQ8/v4zImRcEuj1BWWUlNBzvu7m5KpbW8FeN9rkZUvJBD2JZb1yQF8PHJDelS73S+na9S
ywx+NMAWnfym56ximzZV6bjnOtzhx1ei748s89S4Km/QjNpHMmVWOtPCk/6PbkyvQjxo6NGnpSfc
GF95ZEtwJeBs6YE2Uh281pP/mTf6fJXoQsjHJGFru6iw3F9mM4EgPYSII0N+7q1spUeMmbDj9XK0
00JQoEcDmN/4R4GoADNsHpn0WpkQGjZi2vg1XffzOTxw4YMrclfq91aMikxKTBMv2YumXPXSkG91
PUQ6E5eCR3GuYtcnbSBHrVMaJGSsfdetdLGwy8LcDp/yg6I3LRHLPf7x0gjXj85qcJi7FspkC+ws
3hidGO/BroL8lGkjE15M3YNygyKrVD/iKOES7DRE0vKu40LQC8s7mgHzWxtYWrzuYwiSY/5H2gpe
vg196zr1zsXJjLONRnr4u+J9Mr3j9IMAvHAEMVAuhP7jAxHbwkwG5ceRXFd0l9/PSomSEyczFhaf
nMOcLsqbGozCjN4O/a/8pWbdBDYViEB9Qp+5d7EYGsL/GW4gyQ0dpsfJwyf8JC3dOjNI9Rn1EoY6
GfhW+qS6s1JcpupZPvT99rGYTV+Ydbl1SXbwA6j9cGySXV/cEfTst7TtloMo1d/GJ7pKqtLekfhQ
D1z4vaUg572jN8bn2ycWvf/th1t2MtN+h8LMAxYs3PD0nlINZZYRNGcxao+gGj2JJFb9v+nMhBdw
t3aJ4Jd0E34XqZw0nH5kOenXSrtcDkFXFbOEO5i1PDuMJQoOa70UVuEJIs3Ek8hPwi4/Qs2MwBS9
fAgAv/1MS8tUmI/X34n9VIVlzHRkliQLtKcd7vulySaXGEKVowsRVKgzxe+PH/3mq8o6SdavkZ2q
X/GWf5CI9gCAdyQg11PNucxlxpsNroyn73BVe7UfEKjljs5fFz5IXAg+pYS+aA2hZviKxQrvdiZD
1V+H/LqqtJdiejnoMqFfGVLRGbMuIrIyYy9LWolCyKPq4Hi0Fv4YPwiEC5pXGzbCpiVUpstlmmAu
k8GoXne31ML0S5Ya3USrwh1Dk5bzHumTrr5vtWZPHoYwJgkejEBi6AX6lmh5J+t3I86+nZG1REnP
S6VjilSbyj12deq+75/RU5d1cFAuv4A61YBoyMY1EB86G8LfQgOcBHrULgzLaOzDz3FyOP5eAAuZ
EUf2T+A9Jn+Tpiyfo3n/tYyhom8eivHFmU+cYuwZpxvXYk0ETnhQcGS0Xd+2gR6TgWzR3q4dwen9
3Fkh+qhIAlvhtX/FrvXDSmhzvcNZvOUrllj5ZXyzB0cNnAaIN7BXPPivoDIOJ+m/tLFw/Yp6RhlN
A34LnTiB1TG1cGniILAxUxXDnYD0cEZrgTZVzrzgV6UG6dOunC1NhLKakv7oGENvC2bcqfYmQ1G+
lQ4J/u5tt32ygjnrbH5+sV6e9nAivj+uWCT4K2a4+NbNX8Vyvp6hruzYUywmT2lDvHRadkWenTii
eh/HB2S++5cSpaPcsNYR1DYvWhlFOVw+JPr0CiAOB4aO/u+4UYovmPxQLXqxpDq6PgfAyrWWg3oC
AUTBkbzCXakkEv+MMed6WY3leW92hXD8oOifBDvIocLz+v+TKIvaQ9MNF+racHzuyTZO7dYjFTkG
Jbx8fVWP8B9VnvlODrrydeh7hf+IbjzhdgJHVUxFNZeTB32Uz+oyt4LluqE2lvJiT2tT0B+IaHW0
C8A4DlAYNXyYba72RXEwkHYZ4lqPP++jp8iAlf14epII0A8loSIhP4WyVip1tA6IxcJT+CFa496q
g53Ku9NUIrC8tZ0SfJHZXiPLcSe1fXGAiWg7jxtfxMnGFQ1rqBXO/shIJIORy6/7yi8Vgf8apN4C
DeNCO0rrH/y7+rkIQkjgjqCPuHoc/dTH3ga3CXDgRXf3ENJ6EE2I4DlOjvLYuBZltw50ExN78lxo
+teZnEP/evsKZU9zYejHIFtiinRH/f2Tk11lx62O4FX51D7vRW2AV4vNf2RXX9DNqcMSEq5CzXKH
eemqRO7k2TLnT2e+a9YI8oIdvpHogtVoey4ytGWHphZsHwHZKsZPnws44MPXeMApfktA51AxL5dM
+ODtHAcTZNwxgR1qto+VO2gApC59PD4uPAXPPHmmaA4hLPvMGsmZ7Eny8D+i/v9cSyeUh9Y1gOZl
kJl8ervI9sI6SMt93gQAh7PeJBSJRzSBo1i9Emh0UGeeIPoqxFeIT9cV7sqlvJE9EWiYdRnQPyvB
+F411757NBflHbpNO8X+BLfLApOdW9Joe5sQsZuaGOIfgGGsX7CMNIZqr4uDMopHYE71yw7e+bn0
3LfP7P21GdG1pYJcgZ2E+uS85cN1RZTDARSwTeGV6AwqS2YfREs7t41Sp5/DkmfWA3kvOqzl90mv
Apdp0t9OsobR4vPZnqxroiGH4ktRKTl9GdhEA8F8F+zxRJzOpCbb8bIFpMjaiPAVBLxpBGceCe/D
oUIBvM9M8Zm8O7OSj0rzlrHMoDB337e/KpAxMffLqsJOM6Okts/d7mZhkgRtaFYd9/Tn9+LbPWsk
yM1AffQ7IguGy4MDo/eTGkNCfEvrQzqF0/y9ccZDArD+sLsExzHGnGiay5uw3AY+qrUv6Ak4EImH
VoNf/KSb9tNfpm7WvukgaBcSs+C2nbim7ggDQSpRlErRHBpuqE74k3+seWl8ovNGirjRHw9WrvGB
pUmgPn10XjxamIuoY8vzMf5vd85ku3t87XaGvBc7A6Hg1k2p4LkCPuFmpwODR0Ib8UFgHH3X4vrj
2Vh6P7px1Wl3t+donlRYH00BkOGjFn/yoSSMYhWLM9RgnhnfxDrw+pnJYwlweWPaeHeUue0NMzb8
3U9alVYUBBXMtpyUP2i+eoMCEldjV5fFli7H5TnOC0dF037jLYgt5x3V1jVqcbH6oEJNhYQrNUlG
YcP6KTLja9tZs3PNvb1I6O1j+R0AayF9HugI2i9WJZMbZkgkLImKr+Q7N9XnECpoX3g+1Ipi3CWy
DxstoMf4Ub4Bmeo7/0zSDzRIxnLdT26L0qcoE3tPBvfv2T6gA5QZFriKS2UPUBJq6W/0SZ/L0yze
GkJGETv3ttp0sU6JStz4MD04/xoj+/a2OOFetxxi+pYrSS5GlLkXvdURzwPRgaioBKLzeKZYYT42
bZhIFOiPLZBr3FzZbbl1rJJQLcKSY02XPs+B1N8dVfm+bQb9kpDQLl8LJRauQA8pilUmJ+JA+06Z
cjtiFkblM47af8ewPhUbRNx7KI5ptw9lEp1pNIAecPAK1j4anOExFYeMFOxpld//49JX311+OzrW
ubgrpsEJDfucS7MXAqmjf15WbAKeWm/HVCFb8f6XXX6qebzOLK4MJtZJt/Fzw+qVI+9XXhCvZRXe
tZv/fZ9+f5LbQOOyKfHGgtN/mrpXt0uYye8TKFJNeT5bGj+wg3DyV9IfPQAPwsJOBkNZW4W0QO+W
ys9pU8Tq62jNmRk3sHsnftuvL9X91AAC4zoLopcLf5DfCtpUIdhpUVUZuJAU2XeEzBHMHRrrvITf
lHPfCZepiqiZk1wvoo5MN7jygxSC8rXTuV9wkHvABEGaLAq2D5DU56ggxtmm90sH3luPJ73ND4fW
WpjoJrxy5jCVn2SBDHo9BHRxWb8jRM/NmXSWETT209V8dYDYbUE/wHB6yVozMpsPbG+QbXKx+7/q
D2pkpy/kJ/0e04fbiPOlm/LkQfptsITk659iyXDDv3WhZzcBnf8gr9OsLuJN+2Ljrd2B9zsY4ern
7r75IwiP88QYjtQFn/0fXihjYd4Ha6XLrhJyO1NI5baxTEn708QFn2lAuQGtnoSi3ufES23C1IUW
simQ+CLPFjMRUbKPPJobmzmkmTBVwEmzPLY8PqpObTpxSBcNjDVc793c7uXPynCA5fzJOYt3tgOy
FlOB+TGdIbJvlvU14ids0eCG4y7WoOvzS2Kq7YEEjyC8QXgBK7Dt3E8YSI8iY3fqCidk34Ka74FD
RExgJtaxefaBcshW4FHG9rZ7TTC3ybrhXH+quu/UBiriALcf9TxmTPMkn/cWrkF7Fi2/14owasYy
xomHli7ybi/FkanYwVAcnKWd3gaOtzURfNEPa8wWcIPO7uaOVlFwTarVmYsANSOUkHPDniRhI4Iq
ck8GOt+2XUeLkFZZOLLsNJ8W5g+r9vOyy39ego5ZCjW8utn4jNIZm+hAF22lLIBSz8Ld4WzlYVIY
D6vr7FdJ2Kmz2iop4usBfQK6/JWgkr9BLhDyOm+vhXs7RrL+Xj+n4GQj9CpX1yBqQ2Vm7m72XfxC
9InsXoYpzjOMhfLVToJ6TiR2zid32AvVg/tBsg9wn7MBu2j9wfZEJoG5iqsCMK7JILqFWXvGwHAF
mUpiBP1yMSp8jqqImGssyg+dInjE64QIhJIu/dCeFbyn+iCgPKQD/YmGqx/aJrDMaTEdOMqrCmxE
8181oUI1Tt+mgZ0ZP0KXAufqLzQtn16e0vFBc9SvSYBz6w4QTmhve1A1xEWFDhqbvuutpXiNQUL8
8ASW8qnxcGag4cN8jZbUfCLp32A0PABxJ3NoJrcTwqMO/egBW0sSU+j+MZ15kqHcpuaI5MBu7ZCm
N0or2m7Xmo0MjTABi+e2GYJQ5zS1daGsf7yy2TAMCVsgBrupYWC48vK9kXmoS9VIznCU0Sbywu2c
wi2yV4XYEyW1E7o68NjyYjfNYSHhIxIOrm4u1j88MILhN5aVnClh+ebE+yaJE2W8dk/25XjpddMe
KsqfIvZ2pH6gkrzpwj6dPtyI6CMtTC3jYuylTzq9+IPI1XJCBRgGSnnvLFU9roxsLPy56J9/P2mf
cA4pIHzqhHYcpiZyYrObe1IBbtFPb3myAQYGTamW1mE2qYXguSWTBn+As9K5235exde3pms5iDL/
fRJvQzO4ajfbLCS/8T0DDMHppWQYp7qVdL2WDUmE2bOVRpkMmPnzlALFHKFUxwevzOcAgO3Qq4SZ
o7QzcQjo5imBYvQSpJEVbyKJSkztkenYFryaCzQ/Lc9KRHpRI6F/hCFdeQB2LHOAf+YujKn4PPAC
uyC0sJIm8yR9YxXbQpn5s1nEBbtqRnFlrbcbzCx02NvOI6e6uLuanXieJ/TiIfyz7RRFchYj/sj6
MhJmELkupHulCEymNeCD6alfZcIAIY7S0GfLn2auyRsrwqxQttOlzUHzl3FvE71Xzzy2sOUGgMOT
AM6EOtCOi2cyg46MDjpngoBlICtJJ9m5rlSMY6a5a5DNcJVgXCvYw2oKdRdQwKuJ9YMoCdxN5Ith
G2P2ReNcArQifcxDk8CdsP2DnW6bY9KTq8+FcZPpqHNlQyoBjI2JGCibau9QshtoLn5zm6nywrCe
xpN/pBdl661/wZ48JRC8+WH4V25MtREkgCTZQskd4yLl0nBWJjGHX8bss+NhRQZKOMr0XQzDqzYZ
4hPffrc8uijHfbbk4ZbuaM4h8FSSYdwsDWNeQRuKpgsSsPT+iCPZhhVZwaHkHusfBh/oQwMHGHxk
ubxHOG8VHqjcjfbkB67DPjkYJidV6n5rEvIiXxeM9tqmmRM/U1aKoM0LpKAxb5RARKi3R5C1IfO8
5hZQnfEx/mFOcD8EUFuzYGhzI8Il7AFzC39XrbecBFqcOTxCMegmwOPmxBC0Ww/PTyRYBooXkpse
jpACJwWaTjVOZimhyLlUA8IYPC7LCEMFMspF9i/y2HnBeu9Y/yq/bDNoTkvwwcz4ywLWqh2kx1nF
asSo8znP6LFRcP5HcShR/mhl4knif3nDpMmxcAi3e2+w3EMI62pBaDiaXR28/3muteQ0ksDba3Hn
iX2Qwantr9JqZmwtHtiNpkxsG3gujau7gXOqZg7dhzoIybMnDv8t1tocLWh1C1jLgJJd6vt2AaUx
wPNJY9eRnruxaz8p2PZjglOzasMshTwJ2//xSQEZUX8RvKuTsgbej4nrDG3S5rG0PcIkJmEKxxho
h7gi/dkJqTiMrnz3kSm7QJE04j1aShfH7TsgChErVi6YSY8cf1DoKF5bUStAw8aCJgCD9FmQEyY/
7JxYQX1hp1nfA/8n1dObEG7OXBCbrwuwry38+cFByOJdNiXAgjIv/FERnbAM0riRHYOoczUBMOnC
GXZzB6yHHgZ3iF+7ytkdmFU5mZtkt4RvgOOpnlol5NEjtHmxtqMSO28UMgtxEupIzLnpR/oTSb/u
dC1Dte0CMfIFmmXD6aFlb7NJ1+2pzmxvPQTAfdBcJUgoJ5epoVnNVmjeHQnbH1UOVOcyszgxr3IU
79Dr8TGCMo+WUUZAqmARtQl6FOhovieit0ksQgBrm17adkOuLTokmTzvvguhuuauH1WmGsmWY2HO
/uGFUnT+iWNsBTyhbjuKX/RE+qfWLdVSiz1nMvfj3IKjj6T1TPJ9O4Owwrsx4eQcVrpP1XCI8n3k
BFQGdWmPxdPxhaAL6EYE5w0zEUC6meH85ROKd9S+lcLmN6pQdIeWHPVi4kmvwtHFgfz47TtX3Nnq
b9fB2RYVq1Qtt7KwGVH7HF+h07CgkaKYJ4KG7EEJWsxBRjyb45924PWZnyJHoCOGSBkKKFerm4aa
6oUAggNn4iCB4rRtQmMo5SeuCNXdyCTQdHceogVbFWcLCiJaZak7Z3TpRbN76jN6PM6HggYdQZ73
mDM3Lu25bi/DgqVMYWw2BTji3AL9kz0SHaWmbxJ/4fvWGYAhVUUueWk77q/Wxw6XTIWWnSpoGeja
o+vK0uLvvvRPXtWcwnPRPi6DK3eRl8om9N5biyb3fAj04Z02FX7hUA+OUSKE4b8EeDxsdJfBbxpn
dJeXMMYgBdtHZ10Ww4laIgI8+j1YaeqpGY4w8hhmQeucfx3xuPBeP/EjPbNYfVwvmtuPmKVYFon5
M+yqX4hfTILA/On4ModI1eDFpHw3FTtY1WTJpXI4daszb0Fg1sl3AVsbkHITKjtRJ5xSRnutPM5o
QEZIGcMkD5qQqHZOqFVpBGGbNekaati7JMS8jOIhjABh3rp7PZVMzg01Uoot+p2BSo7eKi18lgMp
ZbmmPXFMp6WepVoij649pbe6Oh+MqgTVY/PTVAK330F1MmfgEiA62fmwRvu1sZ0RNWyU3Q+4o0kI
EK1chak9Ky1t4xl0B1pYq4vJN05lIbsE8FlawYaRTWO7ULSry8xjbUso6bHVYdsswsiARBtdumF9
rCZ2NjF/BVoDxcr3xAc95lr7wmbxYX0jvyCkBuJ4wipzXdFY5OUpvHEblRJCLrVlvstrg1quR3iX
lvmaXPE9ahaZ1NDnyuSU668udRtmZT0ARCVxmCy+HaBH+Hybe2N6m/haeke3OZdxFqeLxMIqLfAD
aF387AZjtYHq1K2RqlVK0ifSna2WNHI4HIrR9CbbNuqdZm6PKs6gMyrMw4HyVArUed8PkpgA+oPL
fJ3oK04ztRZc523Txe0mAzV3b3QjxtxEIsbUJ36e8WnckLjo4cIT5zFtPmVMh6DJchaufSnGl0UU
LUlV57DvK7rR+Lq8Zna8Vd7AYVMNOItKo7ll1e8mzqf+xgwjWWYziCqxlf+S1Ipw6da2EfFk0Fbw
yDRxyt3jQT3vCye8U/dt7z15gijGltTZUofNb+WItR2EJWlLoo0Er7N6XEOEbt4+NhXXt06PNub7
gljpwjFMSheAFIhH9zh7H18kLvNOnhsEeZQFuwhEp0wIV7F0L5ElRvbEq1ZdThMEndCmVGC7HQy5
YXDO082T3i+N4sMn/ptrw/V2BCljhYNNQHESMw5n7+3rM9ymvGle1nMaUqHVKgGBQdahnWB6tkBG
3b1u310N5vhloZ3PIH3elo4b5moEQaH+UIpyZYZLKTbNpuWjEMs0hPDgfGyvJZ58Shj3yvsc1/x4
LGgvrNFNhi3Hw4LqPcox9aeI76jT8GK9rMWbc+7i1tx0nznuI23Fyhl0+iRkTcl6e5qLFJieGbwM
oJb9k5XYscliktppox892OrPwSASBA14ns6IEklJWBPaIpNYwq2HyNFnrxEsKzB7wCfT/mRGPp8z
P68cO9BezHnN7jCZ5+O6MBY4juEHjKbBuVti6jp1saYZSpTHlAn8LSdWAPxI6+WWDCm0wqzZIlMR
EwmG34+dyjaju4wEv4inn4u5AQ03zFv5d88w8uit0DQ591g4tYW/bmqGYY0B6v5NoQIq1pRlJMJ5
I0tDdedvr+slt+BRdK3GMleYE3rUgFQJ1cHmGoJG9cmX6qO/tgDJtLCBIJazhJEtrxFh8lwj/IQ5
nx0+hg9WNfdp/YHx3lGIadjnkmqmkGPRtQvpGxUf9ntcI1FfKxwhgXMbCfLRBcGfNV4Xyz9ym475
D44vVnU5eVtUgJ1GS25Nx0Wdnu/+/e29wyaOmpeiZPzPOWiq6yzoNCwi8UEhqO9M5ts7uxs52knN
WcdpZbgBB33FP6EX98mu5210McvVmDkQ9Jw+ZTE3dIgeqxbLRs4eBjElBNPZf+Rizsas4DsS9+uW
ZI4mBDG/RyuMBYqZCtwvUojEU/90x6GON6d64BQ8m0zuevf473kE+bva0xWE+BC1JwG1Rove65dm
ZI3rr8mVPys9dkN9AdvVvd5AC8XF40ZbsCDA0KxWi1li3g8Gkut39fJM39w22+wQdFqvPoY1jkGb
q/j10lj1bXwvXUjRMzNF5AhXxiEAHCEPXsJkTg51nfEkKN0qaxCAWkDJbuiwgVY8fUp4awPZwl0c
TNK2+ZtlJ7Y8kkXdLlVW5YEbIqmAsQEW2zXdFB3MxUi5Rs073BROBP5aARZlnteFY63D+90TJSXI
DgVnpgHyH62NR0hLloK0dcaccoglJYo5xyb85noLZONfqjPfYo8lnPu0351Zkr0l6CKB2GEANNvj
IXxVtXfGLW+Eh70Oczx5tBUdpvCQaibRyar/dibwWRHIQ5SxyGIN6b/loJ53Q/b6YxVfT6mBLndR
zmaoRrR4p8NRq4mPf2zruAVh/lx+DB3qvSnV6MGNSFymDAQSVBFGbrUCTV9q2ghvNW8bxk+y5GBy
8eYcToW7hQptDK2/lREjGqlhNKBVK2be5LUteGzOAh5VSRE3zQh4JXtG4kZReyO/QzhqbKmj5KTO
1CTMK12PEteTlr9rz2lejg4EO2xt0sDnPJnuNtLZhvwoCIEeGFZjaSR+M8XcW4IQJtH3pSIV2Spa
aRJtm4tcHYMQdAodOx+Qd14KsAlIAqwfg/RLAVlA6DiHZVHOp7M2USpJlHa3EIwQjUwpETthBF7L
rCzqFMV/ba31ZTjUubXeQJOX2g+j6j2lnDjDziGJ4XQPfSzmTFiTuzh+5BNDj7UuElqZg0z53G9Z
sMsvsLFJN+5P3lLfUvN89N4E4QHD+C7SZOrVEWV0bc18XDrGnssbZ2tGbYM1lG0cKp0EmMeQQT1s
I5RZMBMPY+GdBf/9spmNlX+D6RHhC5ZbOTA7P+8/qLec1j4tvrQNKTN0aKn1r+92g9znLBZKksCL
Dk0ca/WBgbQb24p2BldUd4y0e+J7waE7rpPXrrT0M2sfSgjBnUkpPlFtCFx6P3RTlO8CieQHbR87
n1a8EzzxSzATTJqQwsELx33afro9OU+oIKyd4fVI94U0pn66chcSqsc2mfEkCvXYl0eL1plh+xKs
51pI32tML5S26XHX4H/snd1QODnbvBHbWRoS/+Pn6TrKwZICzki31n4J9x+TLS5H0N0K393fkMkp
1dN7aqKUe4maVrDngsoD0fLmPkGYa84UM+NZ9GAc+RCVUhwrREn33Yy0b5Qm/MB56ppA8xrY3dxn
kOb6J3jZvB9UTVa0laNwRM1USA2RiXoaIbZDTyzdUfAnD2rW6kyRQ3oqdJB4Knqz0U/Tey9jkNxi
Uv88U9gs2p7ZQdNMgY7uoX53vWFUIg7pX8pvZi0jwBDKrwXOQ9RcytTIil6cna3N7NnXh756cSdF
puvt3wnTu4wExzI70RklkmgunNwOvxO2fi2G8m2FI7Y2bR7T7SeteIAmyAjJSk/jOL0LWMFPjpzY
oNIbq7qMmJutxaMfcRPsFgvBSndERxjPWsqekHFjKuyogckqCpAP0ZPf5qt4/wEgskebXAFWy19/
LvNZZVTvo67EgoFksAacegPwIIav9KoNFCsmpehx/xJ4fuHSopWqEu4KcbIWLRysLXIr6ynOnNGz
5yBgbNHCtFIKTz7GmJnuvGEj2/KYod7NmYlAiNYLxSV2P8BCrB5JJhZuN/hic1W9p/ufwrSrGRGC
0FGcbbXIhPnm9U0jWwxm9mG98ceQz+3zyXIEI9z24JNddvG3T4vRaMdiYhIfKtOq+Pdijp+fphyP
KbrQ1d/Ip3bLNZ19UjbaGBZ/Xu3+mxko2f5eC8bxBx3aeYtPwfooAe5cWmkLUTSB20JLlUnuz2lF
VtURPA/MhgaujX2b73PL2lqSHi53qUd3nVBvOEg6GAvhM+NGlql0kdqWVC4NPUpHRubWRWNLfvQy
zm/pXySalgM70M64LPQIldsX0Gz+dio4GeBv2a9K3udzAbRVnHXEp24X3TLE+5DRFl8ihN8FMJao
uO8k2WCMTpRngIJJc5LvcYSiA7jmQgGljuHEEqBNfy5xC9TouArUxjnXyr+51ejw09l6qOQGryJD
AQZ9OztLNblt+7KQfeFOSgjiIJ/XKIwTXH3AuLTmz6PTVBtGn66mbQBuwHms94iRi+KICncv2Ii6
sCFd8gEBZDajCpdr0lKeMaajLvOkkZz/uWK9txvTLuGuXKEuHMMtUO0/zsGQNUtorGVa8dfdbO9z
hx7+IUudzwiD6rnfsDCPtjfOn9Hr9ZwfiPpwQXtqymGGf20LTluWy1JV/CswsQq7mZokIin2GdxE
UF/mkDOY6WcAgPnjdMe1FDpzcDdtY3iy+Ne6MiJ8YpbG+MuYaFFY6xqgRpINZgqHI7Tm5XXzlFYN
+e2zT2fAduJeZiB2Tph4qikP+/HOmCLbzBm0ZjaRj6bY/Tat7L5myus6Llawxe7vc51W3+XvH/+o
cTuUXGOy4ro8Ay/ctAfk2t5ZhfGkEujCmE78hM46XZ1W3ku+T+VmKjYAzJKuQskUfEZd02cwNNRe
Cky2l9uZZ3FNAxlDtKTpdyHcwsqyxIXPY+SioVVkaJrnkBcHP6xS9mnrc9nkKHR0OUEXE1aZA43w
hNgJ456mhhTDiw1Jr2RxMSKCS0ObSkRpNQG+8NGAUtyT3Kb/gd5nAvdIDffTb1+PKg3udLAyBrdK
hr7TMnCPAsJm9zKkynI38kUAsvhu6yLTXeVOKvQ0P2dl6zIr004CRxZlttZY9Ut/Tzac906ei+nK
vxJ4J+0sxBWtnOpZaP7VTDfAcTpEmtbSXGLgSaFQA7k6X70NubwW3Dhh/1+RysXGJUDfdPK2MKM1
MKU7vXcIDUA1ulSqXR93gV6jt/EbG1BJuvHaKr45rNJHixJ2Uj2Weosy5awBfsJ7OTVPcWJ4QRjI
yGiY4AGbpk1fbQuDevAW4+Vo6QIAvTIfyj2Gm8b1kLsMcpyPaQHr3RF4d2KFw0PPXdkc7ipG9P9x
+e0mhsheXYWEw6y9m0fHjl9gTR0LKKC/rBlLgGetpFx//X2bHEDx7VOrQMyAvwRWLmg2PngAWhT3
JezC8OE6I8RsrZ9kj4MCPAhHVrUrSb+cmVCQKnDdDtUSiJr/TAnG5bG8WWBVi2NW21XkCHD7ZbrV
VyUwVLw1vhMD5Z3qWFZKXVDYmPpNoUeNu+VTC8LANvvFpwymfv6thDWZ2fKFw3hFYkKe+cyh7Th2
EwNojDBo+5xvAjB8eLh0MwYH5S4a6aUeGpp/k6rXRWFlKLCSjvIcvQjzZPJKDdOtQ8L0hf8F6uzX
SNmL5q8ZtsnZyTOHLy2/V8R7c+MzVCMGuvJXWnb/UdzLKoI2pZ5jbUPR19ospbFGy8h6amCV7ju9
JPyHN7dNglEtaVPmSZVCjl7vHx7PnUNqpVTTSM2hHcZQ/GjhlBJVjsolqCsxcyuQXlWShldbpB4q
RjcRnplBu7zIL5YjRjtdwFceYhvzRuM/Puesr/st9zWHTIL5pFd2Nrssy+VcCPeDDR1UujWJafan
KBXZ1fmiEaxInDO0BSm6WuZc3/trl5IdnZCjAdeucmp6LgCmCl5dazh2ehqMX6ceAQNR2gB970GV
SKU/Tus0qhTW88aImhVGMIJQwBsBzHWZ46h0w4sU5fI4LAVVpx0zLDSL1n9L6+b5H0BD2D3Q4B8V
sXX4E3BnMjWmlI4RzJymI0OoNXchO7SrSAFDIiAay4MFBdOyR3OoEUaPcgSFOh1jiq7qzuHHjAfE
dmPmhz/EXjLmbJITwbTuTDdlzKTyK0eoltMJUzWgVsVfJd5NLCa/jiWtOMvVg8IsvbV1sbmKou2J
OfBEhioVDJ11KZhwpPktPbxIoaHEzoue49bBTbmFee0RZPrgKJ+neGyVoZ78YYicIwPV59TZec/z
9ODAewlMwtC1JphHJJx9MSfH8buz235VXnENC0vyBT9qjMM16gYlxx6WucpXXN2rWKotNUvFEUTj
kb8fL0T06xd9UJeUbQDG2v1V9ejcTxjP8et4DCPpTGIiMgucx63sbHBSKrDTHVFc6uhe45IZnQl6
8ceiAaL9Wf4TKjb2PzY8IAi2kAmaPEsdsLXfSOAEXDbC783G+vWZR/vgfrDNUOoOoUHlt1nw9D/G
EeuTpQSPeiQfltO4q3jgSfmJviC9NBe0FmTQx3HyVjlh7lX+0Wk7o0diadhaOUbuPslw9w0C8LuL
eOddM69pN1b1W+vY7dkzB+OuwZorsbkBEYJcLkwMKY1dV3XLMOJgs7K0BCYe2BHPnAOwLeAX08Es
oMSuexqfhwGxcvJebLvM1gy28Mywvm7WF/jKDB8mhd7kif+deSZnrxvfFHcCbsqPSdApT4MHSSgD
n/P0MzSog6baL1QMbhlghaf8EbqbssIqtcYApWOIBhYSVOu3S1afml3dQGz96EueremyaA1Lo96l
IuN6Y2mXRSjbKavgx7jvnbmmQBAw8SkkEJG1N564ql1oc79j/GcW8FfGWuryLUET0mHValWLuNHC
ROjdb1Op1CNP4nNyL26+XL/nEm9i+RpnbVpB8zAd7YOSTS/xjMBnvwa+3hFWNoioh8bQW/gy7dvM
ahivAJCym/q0GDtSAbbNlD6FI1+2z2d4sZyoDPxqa8sgizK03rIuWfhZ6zICOG4MbSllHLOjGePt
nerN0sg58kee8tgn2nEu2t+8v9sO/eTwT29tre44CJWDJCpDwaQNxRPSfKjajq2Lrk51xzIVHmYh
jd1A5+6zk454TnW02UvMCN+8qtT0EqsBKuMF+EvzotM1rSg6MwmBcrEBUN/+5Oltht5RZSdJRAt0
zJOoux97ujb9q+3Nk/V3ruoQJ6xNxUshEd1YTIsE8qC74Jm3UvfFOsM7wYGi+xf9pReTobwjeNVc
JKhPdrSWcRSKUoe3t9mOVcfXkBFAFiENGUkx0Mdo3flQ+fLwmIr4zhPWv9WG0IWCk/egllU0kqnS
8w04d7ziv55FVYrgythmPFEx0QL3YkqKoI556B3F9gOIxJGRP3ibty/GGOzfTWW4YGJi3jfZF42B
8ZgmatLizxeP5QS2pgfb86pIg1KFGpxeMtTsOUYzL2A+Y8pkYVJ+Wx31TwqojAxo4Mm3inux6sgF
MiNyBLMDAbvz/k6UDNwqAq7ITw2d3ULq/g1HSKNvAl3p+Bll5WJafeZ2oVb5vHhANbmvzBEVVaG+
2uVZ0S4sa+3Vid5AJkTtY5uzdAjrUHPmrRe8O8D5LOm0m/pAbRUAhPSWRXISwvXR9/gGZw5gANJS
JZoDZxXlo6gUbJyPdECNM8wPOHp5eCkgcRcLFaINfUPzB6sOdl7k9EX5BFs3KKu2jv1cao6BshiO
Klew4KWVuVAMynWmZPU1KPqxh/McJSkgYJFNGdYf38OcmkUI1O2e3GmzLtgi5fy16G+BGIq1x15y
rdAn+8osU1NZKvaPQUZxWYqLCoL/80vSw+1W/JWYmCiorDqH+a9/hS10sP60DcKzJEPMXVwjLs8j
favpDd/obnGz7+dsA8jdT+u3gqRrh2abtN7jJDyKt7SjsHZtablBrOYxL6As0qHZ5nq9ySRbnz9B
Cwbehq48yw95vZ3J6DXbWtu66m6f6WCcjpPFpY47zLXse5l05+TKfxISroFxQk0E/KpDaJH+yETB
YfNlOm88PSk51ttE55tWdz7aGJSVxS8ExN/dWtTMT+EO0xTAaASqOEskKfqvZb+sf2RpxJ5P3njT
QezVqGBIKkNP/lCTKoxDNL7cC9+NchZpV9k4ymjmBAgBexGj5E1iKU7gFH855vlxXDjIa3aXZXYO
JtS0TyoVPXVOy7mLxf+CKFBqKSO5HvvS0oOe6DIb9tyek8yQJrCanApxsbfEBk+atHGdhhD7epYh
bkWqOuckSz+/uUlmi8pDsOO5ul/efi+m2vtDVokA5fPLy/7VSmcYtMbu0LGe0HeB8gqBtS+O5ENg
f36Pdqid/vNQ/dUqiQdQ5vY8bwChTap6FyaUXgzdJrOqperAcc8DgtXCUG9xKLWnpmrNK690wwf2
YOut3XFj6d3woqCifNY4XSxke874SZWHU1zqaPb4R3siWxyV3qx+vy8Dglh7NdpjCJ7vMDs5a21e
Oa78QBGViZ6NQwjbH7AkoPfF5iwcHpFivo4kabyi2kXdvWNcb9RiJG3118oNc7oYuiHXtCfl8rKN
xbqxrisGgziplJWWgcZETU16VhW+HBQD+P7/WX3Uigpmz4r3QY2pKH7Lw+iVsKEw5t62lby/oYBq
LOELk6cUungI2PM7cj2qgH2s+87moUbZR8XCWPIH6bBUEX95qHkzmbhk/IGUUSYAQ3G6XgCcmRwT
g6DRxDT23CqUXKez2DvDXo92JTrsF0lJy89f33xKHLa2YqGNJfyU0k2xgAFamjKAXQlQAPH6Jgxs
GYg3ge9SFk+V5pwAvAQP8G5RKc6jzyvuWr/TyXEW/V8zSJlQ4U1p9r/9aLj1KapLu3xAzxkBuZkk
fRsqmc+tS/SD9ocXtUPGoN8UZclZ4jXrEWNmVx5r4owLlTZcwPkPfX253ZtWBUbymY4C/SO7JvPt
vIZmirY+QHRvyw/8F/318AVDTYppwN1ZU2JFtKWalZwChr5Fs1ADOodKOPGgPqiHWuy1wBK7bXA7
8YPFahCyngQIPN4qjqSYu3MD3U2dWVg5w+3OLYBY6/3iUfQs3id+bvTiNIhTvb0GjmZaK73nXQuF
fCL7oR24NxFtk6JCmie5DySVoPXenD8Gf6J/0PIv7mtuK4cSU9UHw4JREJFCGl7wR7hl+6ltcTBv
jMqeWO0jUKtKS0doJwhtFYG2jSA3/P6AQJDN5+Jv1OGxhJUN4g3AGwq50AmV+HAl0Z4UUHIDhnsL
ur3irv0UexO/0Zzr681fEy4I72oWQtyIyICMQApk/MaRcw95U1IdtJkfhUoYzCv7SPEtcbKkXVAc
t1r1aXumoc1xWUM5gg8rzkiqmHNwNxggyfTMenThPEgQrazvvkAB23sbSUbXxWgdavuhgzF45ORH
nRjJ4mR7kyscSFnxcANIWw1fFhzyvEP9ggBDlcimAoQlN6b1EJ4IFBqCwsn2/I+OhajdMTINjfde
d6nYtqst/G2Wp6A4sUVe2lz/JKHLmqEAyThG+5hBnuXCBd4OLrLigt70bXTc9v0cjB7j0oywuf+9
j4h5yqLpiFImD9Bz8bbGs2lz/f4C5+fODHEn5JJcKKfbf4b2J/WDpJnKCI5xfMveh0OHE3cRPTUk
D36g02aEJnxScNzyps9D7WPkkWPaie0bwJCK0qHvbRF9BRW9UYoaGe2h42EyeYvnvfDuuTYDYYSA
gaGTHN2e8ddKtH1XUNOxknypyRaMZbFe88UtY98eMF5eUpWVE2ngoGbLAUeX6ZQi6YRwZtXSml1B
AIaJPwIzaTillX+tEcAbjaGxJOPmxsHPgfVq9zjv4SE8+CmuMtozZOZzTjflXeGeUombMOPf1OSC
PZ8w59syURDKKDaUSYkm/HbnRQD3gL8t3WABU7jgCfO1bykeMgB3oTSgxVtyDSVbtFbPOrEQ+4OC
VZ1c2v6Dw3aXn58pNUFhpNPaF6In1WhTFTfuVg5EyCXr5Xd5pJuMgsmv5LjlnmTIUXZ7iFY8PFxy
z7qkVVdisO/tYwLwVmL3ESE+MXYxKSVRsilOMu0GEauHRiekQPZxOsKbLYeTQnMzQwv6CFYDNfg6
/7CwlayqxpUjwXR4vTwTBmY5wEkdwmBHdwrnWhGQowl6w9mSSwCJe8PhhI8/EQWovOMSUIOAAUTW
qTzSHzsfNVaPjddXZrKvY3VW4OJ2F+C1odelUbuhcdRX8jju1ByiBcr9qgfTO0/gNXs+AjefNgJJ
UjJAJ0s/KSiRGcECvIqltEU2AEwlnF6yrqriabwstLtS8b2CTuTtRZVXKSbCUpg6vkMNZv3ZGFGw
4NMi8Pz0liVyjSfrr5vj5PIZlcDO+5jKI/eRBxxi1v3i4kkPqjcS/6JBEieHM9KbD4ckcALcrAtL
yNiUJLGkgUrc3zhkBMMOOi8ROiMZfcFFD5JgXWfjy9b5UOlLr/oenkqooAxj7lW9LuoXZSPqZE3w
2sdRhHhNeo2AX8rRpSVmxaLzRtAjKRnATrqXl0T7onU/gyEJQ9BOPcuQFf1f9EPS1soKl2ABdfId
e9dR8c9YDKwWG+1xd8ewjUSc6xIbKwbNsKVoJw+z0NiAJLTEdxnw3HiaTAdh0ihjAI3JA3FTODj9
nOEmXAujqDRt6gBNz3I/Z82kM/iRL6v5qHjEl6J7sU9j32HsEtoo0X2zDXWywKiqZ8+9jyzx1x9r
SluGmFB+GRcE0zqqB/ooTeDDZzX3WpWHM12Ho17HDkHFnZswU0qZRGSEE2hfFoFyOGrLaK73ijVd
rJZSzQmnxaJ7vuCwTzxEw7SlUrPUwx7J2jWPwol7wpSCmZa1QmsiI4Mk466dkD40CSO3qGelGSe0
DsHV7pz3B5SlEPE4rB96JJnyV6piBMt1tUF2sHB8rHY0O2rlOn2+6esRQ3H2Ys6VqKw6XKVTePBs
PFBs+h+i6TaQecmwPkZNDVX5z1FVCsv6RutG2rLUF78RmXzv0H2tadaND4PEsnHojR6/KI9foifc
uK7m4rGZQYM3F/6etWM0sMc37cYEXAXecoOaP9pHh06Ttf7+wbElf2wdM7d4QFVfR60gR0hqBCW5
xirVy3VAKY+ZJ8xbVglFfZlf5hAqQxIRBPyNztiuSZxuqNobQGmU9F37gcVvHh55Sm+79WXoWen1
b+PFNPL0OXD676VcvTFOrHfXKVCeSLC/U4kVXdcAnhwQbas0fPaugJXTe5+lLjdDOB6HjBopKo20
9CklLsNN9ZQyluY5r1TGN/C/a+FA2oyIkgHip3sCfRT+y/OLTVW8NQDsJHhsq9tQ7BHIJU9rtWIH
Hbkr66GnuEaJVFx7Phksm8ZTztebOu/M/zfYxb3T+0Bk7YdRRp+gWZMZYQ7TPIeIDnTWaM6RjvBJ
1VE8G8kfpdxJYCAYe/PvKHxy3FRqA2cTyeqS3yQCz3jffGWgH17XT2BWTrZ5PW+Q67y84bNtU5AT
S7H8nzDfUg9PceMH81xifmPcc1B1H3uAaMQkX5+YIp0kj1nxZ4KOormNkaNwDrFshgw64xclv3NC
bLbwc51hwcDWoc9FT/Ia8PPxSO+gYS62XWGCEJX0+cflW42MXr7xkWiK2L2rh6YX3eQGg5FaF6Q2
Xl3H/MXK3K4u5NV8uASfT6QI3FzarzbeJz3K5sQvPT4a8kgkjyIto2HiRrETylOVpNjFv22BgSJV
Zsv2/mgi5mftgnxopyAwnw0sMwRaIwbeI9rOGspH3oRK7Kqf/bHXFGL8HCPj0NCLQVc8HLqBPqW6
WlSSX37ys7nRPsjuEFrdOJtwKDSnqJ9NA5s4cdhphtJK6BXj0S/VDylnxsAUdwQPoCQzcOegrF3L
vGJSl3upPBRi83gsTA+LpiXbm6xm6k9tJCYK/FQAqQTR7hI5lRh1cfTMvjjUXEB2sPNqfoq8SQEy
hJ0VR0tWCahahfgE+v8Gbv0D7pgoBenLn5lX432ezHQTadd2fv+P3xXauoTc5DPJKrq77Nw5rJ8E
tLZLC8ZH24w2a20FRyYaFCxvJKdOOQmnPhDcXBUlcheyhOeVn3iEY1MepG7nw+UT7Z2TGP5PeFyj
jv5usiSZXenlQ0N5Y9s9NPw/EAwmHbOjGk/8HO5QOfWU5WUZSy7oHC9PCPTdCNQMfD50MU5ymVqp
3JHXK/1mv9uDw1OOSpWgJlCuVZSAXbXY/Rm64W7BqVNIswKQgbb09Rs1Bhy1eZoGSoPLruItJiYQ
YueM3xqeyWummDHs1gci4hkyBIgyirtWzIUH0E3cIBFFnradQUF2Ab5MngE5JuaiFl2fXaKV8iUN
ree1+KSHzRR6YrarsUF7xAgy6jetN8jxYa43eOOQ6dKq+bx8Tp0lb8AYXjfakJpzrig9sqW+lnZ+
obuiC02IeJFOuLmQYIGaIpejLJnmdec1BRC1cTp6+z8dC4uduW1AhlSm4njCnV1zaD4frJS7a15r
0V2RtPy8LTvkHk8UgEnyfX8PIMBJvKU+Ii8IfSjEGkyBDxsrEVErIQzjqO2WasFg3KRiCxQwo57B
GS6Y1NP10TaON93rim0eSgywUBcFMsOrBfKiBlFKP78GsjN19ypv5aEjbbVs/qQ4GVnF1WM0mtKl
tuEODCSYsTsHJ5L3YKEaUc7tD/+RgEJecmK/KGRlkWPqJKw1gB9rxuieTrTOLJuKyTInvKY+N1UV
ZndHQvhCLXh3w1XWlTDjAnZgrgUmEMprIY8wNNqGtNSQGrxfbOjwhk+DJztcofKiGTGr/x26iaIG
+MW3v2Zff74q6oFHFoAhy7xrMqVbE4iScxrRte30rwvBrxGJWqr44hRaUU/rnj2psLWzGeqpr9NR
pDwaNjbt2pVm+RoCEDGTosIHDTBmrbqH1ujCG7hz2OkJ87syDYq5yJGiu2lBLhsJqxQmeAASht/3
m/Cg1e5JUxdzYzLZZsEv7QURC8M7URP3yBJ5dgN/sW470MQKS/+/4LD2+BGvA5R4JAF8MqcHxWyb
YQi4ijB/hGHsZ/aMY5trL3dJvt9wRMBkSaimlTJJoMiqofy6U1yp7J2mlnHQuDO3uXDPCQoKtPl5
Zks+SppNj3m06dEybFNLLDiO5Xy3LMvzCv3eYrR/z34vx5mPA31Z+0JsuYHBWwrvu3TZtHR0WWBX
9aXqoGJD8grG36mrYrcN8oSOWly4iXdeaQJj1M6+aEQYECzfhVZhbUkmo3s0Iy0dhyPgelU5e6jj
siOelGrW6DmbxDzhYB6T/wIK+nFJYNs49ZydOGjxCIshFNH593yqKgfRSzhMXiC/3v+0w6ave7hF
wT4SE5QWnQHijL5N9kya2o7Apq3E7QWkT+3ilxMj8fLA0Q9brvlmqaxYM8WTNmXA2VN7ZOR8Wd1j
Poico5HJHQGlDjh9DD5Cu4/8rl5IURNBN6Owe9g2UE7NvGWdOQmAII90bw4e97vBfP2kgjoReYps
XhOjb+rcBNuOVFaPnGWxYGO7SFM4uuzS1sgdZKWJdwhL8cW7sR+aX2PaOemfymOwUKw8YWkj7E3M
9XD/zrY2C2cVurgE5UtMseElcI+TcjiFnK6z/V6VtHSh4C2YwB/xiFi2SnozbO+YPwmv1k9FwrD7
xkZDD6ethiXj+8XkTEq7xrH73xy65KrSx03AhaKASKZ/J1x0ByKLl7qa4TYZJxWtY1rDPQqBXDsL
vD9KW6ssVPk3e9jUsbXuan/8SDQa6xiYi0DhaQ6f/q89GcKOqoUBy47PJ6O/5m2ZJ9m+izCtom8Y
OdtRWLjEEUwM6Osin7saOAYQxvvuhNNWg984ELEAsrUSL4GbAC069HHqiP7UNVPJR0Bp7A386L/O
QQUbPg+6piLFcuL/U+hBiqn+hn4fAoVQ8havXpgBvQrgrVPEfdN4G1Vu2F6k6xLDQtke1DZc7+hM
XTMSCy9eb+qbgCdpR0+nsVIoE1BQ/3VjxZmhozjyZPqwT1wBmZ63EpsBwfLdpj72A5o+Zoy115OV
xqSkPS6FxSBvvoi1eLgJ72EkaBASpiHQY3sXo+bjN7rJjIENRTUk/r4ipqzVYSW+vPCZXgXcAcnh
RxTmeM9JlaBmC+XrxyMKZTlo7xvsdkE/Cj3+agL956Vwxr+rmwFq3AHLAoVZkxAgvYmr2wGkdo7o
Hqo5s+6s3nwT86AVy1Op+QV6oJB/qG5d06lhzb+uIul9KtOE6gHxMSw+4EiLAlZaaQii8A17lZUO
WAFjlqFc6sGyICMGlat0Mwv3ovsM1xDfWnQFAEF/uPwMAV13xZPSEH6C2Dq2mvpIDPkUmDHoGoxJ
TeoRDvMRW9HkiSceGcycUwNCInijo97d3cWayHq63VP3AGlzPtIZnP4kGIMST0FNm5srhCNRoQ4B
iExlM3JTUYc1ZU38uGpzxGaMmmzSosS0iPf0E9vookZ9Adyt5F+1aJVlo0PSdYUeD1xEs8RJfWOW
rrAsKwGhwlpOwtBE7mXNQVoUpi7+UIkPRGGx/EcHL8tAatZPWuYUujf8Q46OwGqOkfeU9ENOXwwk
dj8wpLnEwMqoROCEVSwguF/XPGcpoPn6obTqYae9tPYIgpJkuDU7Qe/6orqbdXUO7cnSLXsv7h3n
yHWKTcdNVqcJdFK4JwW8WTthIzr3gCntJU6tZYMkCWxxtFpbOpgNx0upQD1LdE191t8bSN+QAy5Q
6hIxt3tZqsvPwZH6USkfkeRN3z+56ViNpaMQ/BcyklpoSGCjb3B9TjuphC6QZglzLdXRILEJHcOv
nOrj1h4/ks7frwzomdr9zRXxkaM5R8EO3AnA1nrhd+s5HHPNX8FyIPfQVelLkOQXnJHADmN+r5Gx
Y9rLpPiRkEY1TGaYm04il5qcRuZzcagMXVvAxbE91C1gVjZ5sXTgrCJhXghMhgOn4TCNW1jeuHkD
MoYXUWlmcSTfJin/WA9snXQpuuBdw7z8Wa/yLzCsp6ExKrtjaNu13DyISLk+ac+BO08WRLzNq4a0
W+++x01Jm6zSsYdUudpG4SkOyGV1pY6NFqfiZYeFzCxHcPaGDmXRdlAHXzMJ0t9dg34RNohistKJ
4goUv0piHdY6zSmZunaw6yeVzAJV57tF9whW7UbLA84+2JMBhDHqSIkfeWqPZtbsnDtFLNeNe2fC
eHcEpCjiCzx5ZuvP9+rZhkoCM0P0Y5ayDnj8WuFKsH0OPzOgYW9jJS7cHdr2Drf6v/UjN2Yn07k7
izGSJU23bo7+VwqaK0aq4H801P5NBriFELhX3ka+vdjXIIHic0Dq0QffDHqf01nbTNua9LkPgWiz
MXYtljwtFxhuCFFTvekF8+pcLfIalTAT0wxHLSd5aRi+Rr1IIt/ol+KorNXr6B3IKkF5ufW0dSVO
G3r2jnXJo/h6Nk5pQ115/SgdOSW0783WboYd4cjDIuM2yv7h+4AGs6tLblhfYgZneqt/rINZSZCg
puuU4p1j8wg/AZdXtQSRaaunL5L9ZCVcZakFwMISVjHNLOEEFpHGx6ht6iwJSj1NXXDxbSpSk7GO
211cSRmCk/yYO3KMtZK6Muf8UE6sywQ3l3K3eF1DjlIIh66jEvQzsE8ux/J6YozgxoboeZu+oG/w
okAUUVeeS+R6JpqcWCjVrul9Fa9KVH9L2+4qoeT3WzZp0NhQdmseyztGTwzNo38r36LU1FGbs1WO
bIZVYrn0/rx7zrA9cS5fqKjFaUtqu3xWFaGtoDc2dTSlV10lwVI8hKpeyZ+vTpEC2ba9H48LPzxP
AxqiMDI3XGNMhQMosz9GJk/46hfTUynMOTZ3uxKnz8B8OS871PMAsEtuNAi740/f5/vMpUx9yxSO
226/ts9ue8eno5WfPM1orE5L2WFbWqF/56UrurkCTUNERba/ZO/oLK2892tuOr2YUTSl0eJrw6ms
B7RlcSqzGhyPytV0z9fSNfN4SHILLoyIp3Sa3HmVBSMFtMYKfNGMjU71zdIURCAQEHVOHKRsiZv1
dEyplN/knIa4ANNjCWQEDkF8Bo/RZ/mm6Ix5sLk2xF3Awr89VJ11KdjqUfsYK5U7v4+kijX8srV3
H018fNKmUHzKDO3t8IQXe18AjTF1d7LuWxLKWRVlqba3i7sj2zukKiX7CNA/Ykl/AjrOcisTazUh
gOiDDlDTH2ieAp7gvqeCwcEemKZ1yV5D5ONctuXEvCmxyD1+BHc5FHIZCRYapN8qgMxUOmPtQiCj
+XU9x8WJmz2TOMV/1rZlUGGDp1jtiL6YuJVj2sqJhB3EOOsnav63G3KL9nIaFbLupr+lBuyJUa2d
dU44wtM04aJAbAv3lNR2IVcIS5SP2XxoyyM64LI5ESUj1FQg1CGBjnmIfTQ+fMEqZY2XGP6epnbP
6F9Vyu8+g9XyKIyiFsKryONkDj4CXgdKlbQ2OORLwMhATcjSLyklR083J3qP8R1BqYnQe2KXO366
MKnofZMEMdyDdSdvfKgvdMP84m2X8YtYPy08QYc/Wm8NMjqhUI/leUw6FKB+KwCM8+3/txnit5DM
WSefbQuF4Ztntw/SSmcyT/4PHO1Snd/kXhRhS43j3PS07axDXWLZzWhFaJqL8e6rqrcnENbmUkJS
MS0gBr55niUcneNxs+JEf4VXEi9m8iM8xlkMVpLPuNDsqbLXkjYvu8a/4WLMTnYOGdrNwduY2oyX
kO0qtMMUNcQ8RpSmrbJAOHVU+DrrrLCi1GSOBLRPutGjz3fsyF0Y4l2Hpt69Ar7TSwWXZZx4hZK6
hh9WbDKpAlow0SELxUvIUacN8+fLLmLHWRTb/c7dP/DeIO+kxdeAGBrrIHAJGt0IrAuVBcz+o5da
Sz6Dg+Yi80UC2lxxkwP12JrfUTviJ+LcubUA23IpjiCLrG/r89WmSLKOUHgaGB90i66D/G+2/TDN
QKbFsjW0t7vWNS6DNwk0voXqENkTeOzs+/SfsrfozmJFoIzhXQJxF66GrMQw2yAxtil0ykRk/pl3
BLqONv+X4+Y9gsr6I+TIIB4O48PQ1lMdEwOe24J0FXv8IQQG82MW8RTka0gyeMn45HCYoHxS57j6
D3bmJqo7Fx1NynV+cYLw2/uiinzVJ8hyXwLQwWURwRHpr0P0qs7qRAwVV6G1sGhY+mcvumej98Bj
Q8wfboMwx7TUWfB1wOeLhDjCLwDdwFXr4Zjdfk4fRl4lP7F+sGFjBFvEl9UnunWr0UPRefcaKhkW
UQaA4YjXUvlwMDKjtESywjhieh/7hjnkL8We/0u0NU+m1bm7x1kXO4Tb+mpoFwtAYepu/rd696Zq
iJFjdsswdEDxz8PmwfQUQW2/jkSgE20/+TO1aIUqxUCV04RpZqMRRTRb0cEf2RXJbk73HEClajaJ
gfwHASuEZ8iXHooSd5p2EFtAS5lttpHqnV6Rf4mlcXCytclzcFmBX9OJO+m1b0p8fc4ZspBjlj3k
Hro4t01572+xV21Jo5UYUdAlFOEc6q4VJ+x8o5WZoc6+JX6cJh8RcnA3as1YWp6Cj+grqIIpe2ps
3cE2JXSbLYTSQdDlQQx5LtjST8rVQvH+fQAUaq6X5xhnfOxbBKoJZ9yV2imbHCJcfv947jOQlama
yT9RsuTN/db5AlaFThDzq6NmWqWdhdzeN4f/mvTF3i5VFz7do5Mcwx+YErifiOZft8xbCqzvpura
vLT2RMlTJkgoaYI31CMk9wVdIGJYSEEDV26FbbKzsiuWZNinFFYXNEX41LeDB8+ApOv7QM8HlGcT
SnM00NKzCDu01fuZzmZ8tkLEkqEmcqYWT0sHe4GHE0R/oRPZEvaWhbGDlRD6d6/EFK1nQV+asNoe
HDrWoop4fJK7mjjyHIhG3gLS4P60v3xW4gYl9tRtrooz4aNPt/OSuSjuq3Q1JH0dXVn60fenS/DJ
sw9O6G0PHgFNbNU3dA7uBc3pKH9eNolOJi5hflpw5S4l+HTI3dG6OgGBspwHcnpPYHoyPmw/WDGb
Wh8VfH/o4XZRznlWXYOZ3Li+hZI865bRI+DL1I83slUJmcmAxjaVPcJSL34DAsTKQEWRY5W3X6kW
79WQieFkRhC9ArD+9WjNRzbn7oU11FSxNTMWK6yZnNAe+m1yz2zi/24U4jyRJgBalo9d2yrgRg0G
JTDmSty0drUbqOcl3/E98DexHKZBzaLJdH73MtE/LAMGs2UPbZDKnQppFCjL/6MOIjQSeMIZsaqq
SpfgIjf7OMPhwQSKSN+9xTkB9t/kWP+uiDPz6hFqefMpHSKhDgGX6Vz2K12hlSQjdqEjFsFKA4wO
7Ib+b7l/8tBQJyrNrDQ7gRXdvWSenFT6TlNa0UAWq9G06RhTc6EUqr/UEBNZNn4WklOGT8dEwTj6
h9PiF4VXavlTBcETO1jKsNHcM437I+S0Jv/YQKZu5jCKdkFSxOo4rOV2rWYs0MgfBywiYCB2hKC4
hcyFxBX1GgsF4UZPY0+XOx3bTziaC4X4ofTmck0CLWqMt6kBe4HNbNgctNPZNjOhatOLsNBdkc2F
RuJ577iOPhW5LUMBXWthgDxeXXoUtRX+BwkQOmnwX3wGNl+bxsZ/fI/r0YVsBLL1n5QUYj2Lfsk0
D9jEge28HjwEUpcWKeF5I5RqdyznINZaQbfZG0STGoXezwNcQ23oAuAFE5eVa+D7AvfbF+7NCtsg
Zmb/ab3kco/eAm6UjZ18im476oXzPtlj5dGy23eb2whvBcyS5Hi+PaZ9nnVhBr6dYqbz0VkjmeSq
MSkHuA4HyYsxXZ44U9eKEQFgVsGW2drhekWs4gzB3Bm/d7r2LbFJJ336fTd08eNyMumZdfgwVRNF
/55ncmbBZlZwcnrwKIQ54dW4nzkf5/ADmEebErcMx+8JENBmKZ5QV1QIQArETSzhfge/FBHT6Liv
KRfxe9jMmSl/ivxnSR38S3nPFfpyodK4F5AsBAUVO0XKCN9eoigZpcNYme9QsRv4PZ32u4iHVonY
u/oYyNYTzz/oCsZNwA8W5zckFMOOndDCh6Sb+L6tRtZjwqWo7KtPwQVh731B/63EXY5CLgdz7M9t
ckGODnHvAmqbjbgt+eH5nc2UMjUOmwovsh3cAsWQleAoclnOYKhXKCuqR3D62nAzsU9gU5aM1UU2
Kv8TyGGrwDcgjhpfS82Ye5vQEs/lcDZg9hklpLvAVRE/ujGLzr/XdyRtBK0AmCnpV7K/gGyzEv6u
+GAfGwPOVwuFwXB8DuVVO20Nur8L4D794q/PLgZG8qqWXtydrFy7yBgrkWypBVgm9N0iIIa1kXKH
ZHf14XOyN43lRVnnC6lS7U4/trFjnueLjavBORBYJQRodIemvJ//nBiUD45TH6PWsigYAsfYbJnq
YClXOfN8hukZXWSPGaf0mQEUvnrp0z+pE3xemZxEkA1UMKID6XALoZi3SbrJqE/pZVXaQALTBTjP
2NG5wmDmbV9WOvtebL9hkJw5WEFsyfqTC/2mlh6rUVrS2WDTtbFz7ZHK+da1N5hJ07+JGYACHLbr
LSY28Fs5A0vSf9yZcW9q2luCXQJwZ5XXs0o4ieZAMNW/lHy4BmST5nD7NjoLSMDsqc9Wr5dk1EBD
ENPpuqztF5teCa/IaDS4wijl4l8bhGhs7sjIY6rDWCiMGksxDWaOjiCi3WC2vwAV9/cWHg4AmLLi
fxUTNOMVyJ7Tt2bv+0LHG1osJZWXVHhHZ68EOC9KDRaNWdQX2a8DHmks5UWKAbxasZNwv1+Ko5WS
dhF/NG3eoOLJu1lkiUImTj7ewkm8fAt26TJqiXfErd8IemfO6XsfXw+bddA/G2vshtEh9hWZMv/U
gO6hL9fOFFyzDQxrVPXVikRc4DAo09JeGm5FwwUXACltafjN1f/jEDI5MOZF9JyIzjuzbhMdwx8b
KxwF1mAk3lWAHw0ljG43vneczo9e0sx4BJCz7iwCdwCTGEqKN/pR1UHAt6KX+Kg1QwDYKoFWXrKV
rUXx364GmKSCe1Zky/K9JVBEcTkrDBZYRqLzROYF06LQgKMD7BcU/5slyy/nJ+qpPIi/LlmxlwT2
aMhJ/SNkqkR59QozOwilwGnidazqb90tjdxDUOtkBGeC1Sgd1RBDKttZVO/HAc6Ha/bXpyj8CDAw
KZKbtpREH5hBlFpgPZPuLDCnERH7lcz3fDYzBeRsrg64ADkRpewtKWuWlAbsZkGj/tIqjpDfWYiS
5fUKsNAvjjEesKWv5JvOIILKzHPIgvEJwBboIQNfcz76X137csdvMHi5bpnjOkZe1jEMq0L1RfII
LUnjlxEd7sYoc5hYK8Xm6bTfz4bYBRaJKEXFSJ3biWy6+gnn6omPOFnvcz+8On/hEEa9dPnLiN/p
SUOVvyN09UkhHAbZ7ajA783Px7cVCOMKXN6djiaBlFZk33PPw2XcfDmQyuB20QEhrwMY60h9yKjw
+8xaJNlOk0i+8QoR8ALu92bmLiWDgFnsEAf1aBoV4Txw18tbwPG3HW3O/VCQLjRdkudL0gc9m7TP
b/cU8SL3i/t0JYFIvv8DZ6JPzEabJ4U86rKm33F+UfSHSetqHfPOd8L9bYti/bmUpBTNdk1UdRjD
/qVMyQQ3Pq3qxxhbCHC7cIhU/CLxdzF3CcT+yIBDRX3P6HMob+T0FrsDwZGpR78DwMiQ8Kems3cc
vh7CFW0i4yhXUW1e072DQ4Hq5y+3u+2M9kyB2ySPR7RcHES1b8p+GVHf/BpKD+DZXjzRuhoxVW+9
L01oJdpZ4r4PN0L7yD05mlumo7/dGodVpas3yhB4wimaLnDN7ZK4pjhoXXZ/1r6vhlAYe+Si7bhQ
pyymQmSENfZ5BMB28dITeOaMOqp1kb8NwnNDumMv4UiMm9dZc7yQWemzyNpssY+B0dUuOvjHArNj
d9jacMjh5dSebshZe0pdhESPsvoj831O38Uo4vfGp+0zC3ChiS2lRjQR4MiO84V8RhCm3zhIMU/o
QhvaNyZNjujYs9dV51x3tNqykDXQxmCE7s+r+pXgbN2bg8YyHsZb3Z1Nz5CN4BR2jMNqUGMgHS3D
wqXe1lrmLO6CK8YkUc6aGDtiw0Vk52GFpNRBpTcW5tJy6HYL8JXleYbsVR1YKWnkHvBZQScB/XCa
2U5BAee15HJGKduAUbsIiNy6laUE8VQ9zjfFMUNs2HUNnoMLQjumXmNEiZ/Q2pfV91T6cOrm5OHw
9RIb2MF5o4H4tNG8sNdDVFnnboOruHcRZQnZiiBFUoAaOKGm2crAm2F8KMN0FkSwiVwWjUiuVIDD
ciC+kVL/gwKZWTfHR9d+7+aHf7cmJDkY0WIRois+SEa/HoalypjYNFzEjaxqlLjHeFb5r02Z/VV1
fnihop0fys8WwdeVeuYvyDKF3KDapFn4RbQxAAFc8v6afx8iIDTxDz5kwcK1kG3KksITfGAZTWWy
sXh7lZolh6VS+V65LdggQ2nHRc2iSwEM9t4AyxVmjP5BHsNd2cWKdz03GFLG3QOJvw7Q3MsQv87P
/KJCNzss31Tbe50b0yhA6/ERCkSVx3NcY75HpsnC864d1TSKBbRexPZtmuW6YoQ/LU/A1TPzk64X
DlqWteWqu9DrsL0hhfxNC4IZSm4nc17w44FQBK+i5yo6qoc0Y42cm1IUXOKqwM2tSr7sgEYHhNdr
XTAf9MV5eweuFYG7auIyEqmhdJVzfzoIqgrk+oHxdagRyLa6l5ETHRUZ9nq2ul8NLwQZBdPyPxma
ZpPo1ptFvBjphirds/rslRA+r+zGUAaY6ZCCYvFaqkHJVLM4CuAPmihlhF++ZWMjWOGOoI6OOAok
y1c4/koR4OF7nRHkh/8k4aeiuP4Fv4mdZSQw3MExo4YiXyOy3sbRT8Gbk8pbQCcpB5uH99Ge8QHk
ZQ2+PpdHNnmVImlcQK7wC2tj4gk2Z/3whoVE/qDUBk9zmYGVuAgUNEgJldfxCogwd/pxq9i6UB+a
wk9wDaZ9jWqwMVgK2BPuUHDyadOPzhz6LYDp+1RlzvnBXVkDPN+xRFISH/k9YU902HWIyEpCiXcS
yisMmWXGGTwaX3k3KW+nbmgLFjMg+bO2o8AdxYwow3IB4bUAw2jTaFSUFE5NbXuGJg5QlJhgnDcz
keMgwHvbDf54cI9APTMQyT70eiG2LwwuLPitgRaz/Pz0roFce3sNx1SPdmPg2oNRM6wryCUR9iMJ
A0fwW9kQJlJegG2mwPenwZ75qFCPnxGU2JAtkZbgELedmemKrQ2CLdlXSQQMgZZe/TroxrFHKG4U
qSfJjU4YAFzJ0/lYWjf65obIQXDZUBN7zxgcw4zcszzgBh2bPBBfm4evaCKoN1tGYXbA+nSfEoA1
O1QCcRvsP/yHVleHcFyvodgDgrRkdOxMHnKkKRm6O9vZA+trmrl9+xjXE1XiQ0HrmtqvO5xzrDJX
8jCnofuqd4ZTbB7oq6mTV5VuRqeNLRbdexn/Jzy0uTyjH0Lm5Vih++qr/J3afHLZW0HhislBcQdW
GYVZw3pygAiIZc0R9VHcOPKbAGO563cNoYAHg75zIpp0tTOWa/M/8DzqcPXQTprKaNtUCRFruv41
2Iip4trkoY/Zlh7ErNq4pPXuFWXJyNbXSNHA2y2a8b3Nr+dSXY9JmXkWmYR9Y5wJFvlAoipAkzn3
VVUjevNRibgUJUCD8mDsJZbISrnEQwyBocFgwR1osgIvIJ3fyVzoU2R3m06EAgdBT+55B3RCaH0i
2h2pu8tT6m/D20kfILUhI0gWf6kZASC31j0/dBlnKRaTHeCqXGtJUAm7/8IqrL7nzX+dLySYBZGI
am9No+wOBQf/EDj2BIbhtLTUQNwZiUW2XKM+5XyWv9GPNnhtkbcS5y5EgnUFhg4Up1So4NRfaCBA
NmhXIYjkzg+wwKfsoo6eHnTrDgrxGlVwRtCDjjD+jNyZ7prszBjDT0V0ZM458gnk5zsU0praqx5n
ERtsNpl+2maN+dKiAQpDLVYzzg21Lnmb+Ks4495olkZLJiSrqccMMYSnVBAw7+VOHWXq7aLeL0rd
pJ2HqKVFWNe+sZGwffzNiJ1AjHmPfzOo+OhIXswXY/MH4mR4C2Wzuc9ZlQfRMVwybmZqhqgFgfMy
iIvoDO+kUrkFMreOo8ia8/29BVHhC5qFWpdNbPFcOETGITBCefRQvjWogD3MWWwSqvDhj9Mgeywf
I7RRay7VCxwSoIqZ19Q3j8XHYRXyWloWpoACeDOn8CeqjL8xbL9eMHWFKnYof5sMUaxQy+rQuf3o
3jGhWBf4k3kWKiPeUaHyFnEG7eD97e/XMAsBNczdJ84dtWpjCe2Jmk5B4VfJCuaktVDKMpmRYl3x
L1sNjTUayeAFdU/BPWiHfAAZjFMzIWS5G82fj1/lBTau3+WYCEazH/wjaPX+LV9/YSE9VHTfEIXL
x2Sio2hlyrVYSY3GA3M7lP/SzLxslrgCbVGiCjFvt4uD6F8SpKGsDeA5c3zb/x7AwTSnuLfhLZyT
1Cd5Qi7vdYTXXeX8+mvzJiGjqx2H8nAoX0rObXoTTnXoiCuGtcUjYI9AFJVqkSxy1AcQ0lUU63+v
DK5+i/Mxe6eA+wMObJYAFFn6i6xQcC/WDO3GMrddVa7nw2qvQkvqy/GA7kFZVeGfEHV2hcwHnPAM
Y4OiSkFqmWFxOxaziQDrOniJyigS5WFHABFzl7fXyFOmfqV4p2vfTprIO+qBBI1JK5CNEBq9Jth2
k4e/O7g4wuGFtbcyJ1eBZejg5dCJmaDyfiIV5Tif5QM5oPqpS+U1REjvi+DtjgQDS1vQJghz4xmU
hdcPGLfOZ90uRdEd9Pxmau1wYGxIZ11Jhvi4r00rjbUySIfPuSJJxBtWIQlm0z30bltTiUB2Adan
AqsSWB9tm7G6927Ve/YvLa/QTJEqpZjzvrTdZiTsKCQ+0qjGPwhkvdgOGsJuP/SFReyGBEcMmwrV
kO/rY4Ffrih4Hgh2RQ8XwuVlRfvvHySmStvCyBW7Jlep59qb5V1um7GDd1jaS58On004I3dK28xE
mwjx8XtE1+ypR/jgRNrT7BJL97dWd/2D6iWURnu7fHqJi5oKdmv7XuwH+3di5ICa/Ci4n6Vkfdlv
Aepwem/lDz/VWcjKAzd1A9hYK6sjzg+DmHxWqblfXobBfhZTXjiXdbdF++uxiPL8oR5eauwwpOLr
myNvrM2TKImurl1+VZvYdXLc70z9NdIScKAKo0Zu5nzLURumrlFDirakbgAe4xL2ovI8ms4p1W2Z
8tBFnWvPmkazPMpVndtrCDRiq/i2BXm20z6Nf07Mdkykzm1EVQADL1WXyYX/XtF/5Ded+fCpanvt
r94/sjXF5fyg49vDBwCTpYGLDhtI2YDSnxBP0YERdJ2VCP0Ce8UPetE4EUYuYJNhcaER7OF+6oUu
7uiqIZQpeX9N6o191wqx8i/z2sQaOzfdIN5Y0hvpWEfnP6C8ym47Not9mHrdY8zBQriwApC2AWYL
Md9f3KLt0UGYvKUZW1J8KKQcRS6eTxjrIZQAwohjE1YFTvrXCtVc/6K6RRJ5sbYKy+islgQPIB8K
0Xva2XVDne3WLBCp/znE4qhdW7YermDnXvk1iwikvjS7hOc1OyYiV8lCnn3CWAvRzEHl+whWfROp
j0EiOi3w9jeVL4oz3fts2TXHio9xF/lHtuE2C71/GocfyfXnZgDDSaNZpVpnVQzsiXK8LKD0tWdD
jsFsAZSRfNWte5/N2HSICZNovP0xs4iClTtEdzUGksauAnxdInKk3pM4DZOVK9sNSPHjzJJjJNlg
0R0XPHKEeUAB/zuhUi0cX9tLmWGCD0KAnmUNSOijA46kSd9Aw4XaFMtJ9g8AiH65GQo1PFuXzDBR
f4mPQTOClujEbAeK6TQElg7sfEPCI6oHU0eVKHn2jeveKAAVBqm2Ov2cFBvE26czvMRogqnkCnx4
UemqHK/MwJhB35AbMelnGjeP09s7W8pk4dLJT9OXx2+QGMRJP5cBmx31OlSZQfMbrjTavgiTxpl6
NgNjtgTi203KLmWkl6DpiU3JH8AL0/ExRNWBf522ARVHjQzch9cBPvrdcrh9zYMtpEs/vxU9lLKs
aeDj9SfdGyq9tz1y4TDHJNj3N91LQBcp8DT+FGd/lJt/JjAw5YuZalFJoBdpEHeNhOczgqOQmJMK
xoMPrSqlmEi5C6HkUrtzgmFsG36aTMTLWWUSNgZl3VfLtG5Dto/Iw0DBwZMk6rDlMIJLwuaUIzie
GQlzCJqblyFFZLSTKLDzXhfFdu5G5bm3Fy8vF7W0fxrCCP3OMTxs4v2mi5Xee0YRKdaOegNXro0t
sZ/Xm/SnRSv+f9gp9TirPRABymiS/+c2PmaiKB8fngyuEIvl1I4QdRLziYJLo6MiKXXQVNzWWRfq
SrKsoEpRwYXS77Vbash6BXiUmFOukujWDrmRxQ5I2JapJcLpLpQ+MbMm4mfunXv4iIj6GcjVMZcr
QRe7vPgJ5BITQuCFNZGGmAP/raMfWMm6iCSu6G+sGtIvqgVmoVZWoSN2FuaMsd/zL4PnAMrAbM8E
w++Aew3ojPjjHJswXFfAATEzfLESJrvaZS5G7T1kQfJ+BFwXmgYlylQlBcAL1onGQxLwHY6OD1ad
rbqj47cBMsTNGvOHtl61m86udYEKKXEcROIjylDVyRXnIpw9y50HO8wcBVErGVcHovLaRbS/qNY0
t1xCS6ZSROePC200MX+ohX2qE1aoPYh2YIYpmu6F3oa/W92/0YfY/FZnsq5Avz9N4G7EWViLedMd
cZVDg2kQOJ6kRofbsu+g0XJ0CILSRJ6vyTHMGJhaqvFuyRmVz4NAqj2tt410zW0uS4xhfDEiDJBH
PuLhvIEJZszHZMpTsry6ITNuLQ0lyr3u1NOclez5ABE7VKaZmCR7U6+uEpQsJhbqHdvKhQLvoCPJ
FyNtwYB6N3J1VX51VG7J7tW3TQi3xsKkTki+X3ks1M9cqXJb1B1mo5ir7M+yjrom3NwjxfhPqPF7
F6Mc5il0FP/JPNHI9NYs+kuCyT4ZKra23fQGP9e+wCJBZElhd1SEQ0GfF7lOjKvaOIRHT0xdFEmK
KRH+UmhsKBrPaJO79Qr0nu/sCABUGqSHPHvF3ODC252y+FvhLwA+FD4r2a0hMILWbeM5tTomAp0h
vyqmpjNRFjyefD0+kf95OMkxq6vBFUbIEkZ5KsGviqZsAbVGQZZ5/oO8oAl9tl817rx0wjKZu/ki
vStIeWHHGuTZPSGMiM6qyI+txkVOFEayHCACDdgQjJTe964sAwsER0098quTBliUdcz4B4tl3iB/
ipg8Q1sdRVhuSQ8aDQBk8vTEQywaZMU+r8QmfVHDuH9fUU8jJpce6NAYg8M6h+68UHBFeCpaPnpZ
CFqhTCjz6eIJScTzxJfc1Xrm/+D9Cs3pbbf2wmhMDZYHLxa0wbikxdDnQgP7FSMLUc7ROLjvS45T
t2rbUnrV8p1l2OC9AH4LXYcMlcAo14OGdPY7E9l5j5vlQ2kmCoUZID4k/9t46ZZmTJJJj0fNoqXT
h/lRh+Y8T/e0M6X3KUOCngGDmA/KaySd472xvFEXBZHddnSz2R4OJpCxPWc9hZxSu2EZjpJLn2BX
fgX3YW7G8UJMw/GQBGflN7fpNCnP0/X1HAJaoLmtEpKEO4Ne7ckvAAcFm4BeJvABB+IZh/+5Fvmz
0INbYN7jaMc712hIgusGHzx2z1pwGWLcE6+5WBbRF8GP7W8iIR7fpRPcENxKugkSvx7qR5lCH7nl
l9VB6SwTalQ46mV2JwbIe0+GVQP98jLxMil0amWnmONCi6aAwMLwfKmIiRvoQ8bex0N97oUuuPfH
VLNfMER5rKcwH2BCr1dQXF532orwirRS9SYtqZKSrbd4xaSvX2HjYpsI3QimBPkXu0yb+39J0OeG
Z91dX5hU8s1Y0M9+A//eQYYUHB3OJBIUvWXfyJzKvzoJVFlR0OaU2VAnWHZdw62DBDv3jjwjqDxj
V0imJkodoUc8lisZ4Mi5CAYuPP5PVMqF71+wqAlmbdMIP3TT2fUzi6eK0sftoX4tPFJ+WsJBDvYX
ybju2QW5kTc8F1m8uzwYYy1nIYKTNfPNiVE8kOoBgcPYge6OqRDFJy4LnzMvyvVdZN0S8KYyyKiS
hcg82k/K6vbS4A96Ttv8SNNelA5d4eqvxOu7xlSFiiH2IckqYkgO8qPtRPk3PsgaVch5EG4ks9cS
9esmHkgGi7MunUeyOIbMuwtXxAoLJFPyeRtZzC65hZMo08bZMuf8ENxeGTaT5NaFKlHW/+R/IJM2
/IEBOdDcS384MlqGUCzIPPohOXS04B8BEguw+qPAecSRdUzCMyMW4Fws/yUQTpW/5/UgAIJ6X1TA
P9RWEAjr+ayluJoAbJ/zvcvIcs/QDj4uHTlwcOwNJ/Clf6PM8+01K7wzoC6Yd0HDN7VtqJJKpLd8
OAgLgIGfMpcRZ+v+KFOzOtFot1TaGb0wwZP90Xzi8on2ECecczUzkqrB1GVCjaeRUSa3aPM8nelH
HU/e7zPQTMq0sGzR6QiVGCNFeSWYajjRoWPIjbz6yGz/Od/V3l/zS1VUeV9lZ0DrPvTvzAj+1w8H
9Ecel4/OcjNKO4uQbmf8X73HRKgx4wMr50+EPzYpLKcrv3bZOs2LDZRBzFCsSwpih8sTgPor+yP3
cugPOAhAk0BN7DKg/zy3HHDYl/zEF7gxwligkUY9Sd7O1JhelM/mQ14+GQvjcbY+Tl4vOXftO18T
wqrLO4XCNdM0k+2lBmDeegSCZQtPq0kE9h9z6wGvG+5aboSr/qnAPGQcKaEfR+hpvlSXWIF1sXAL
Nk6DZonFtahSuu/8xAklp95DBHIsXhSJn8ePb6qc+2sEPw/eIXA95V6M98elu+T7L8+r6oF0fKtR
VCliY9z1oRvN9LobNjP8Rc7du8myJIN85aANBXhtCvnF80qxkI/hskmy36uMtKiLB8MBQBoEURFm
sB9HvtLiF3NAqjtQt8Qw0veYe1YwoDmLVxxCvDAfsD21JYTSdP2ojpPO+pH2AVAkd7V0hiBYEeG+
qVfaMSYH3+9JCa55nUWt/BeT7mnoPIgEQpIgG6QAaMif06lreS5ChFkbxd5yg9P1hxtZM7xkHnTU
hWaBlT32ikIWXkKrdrlM7H5oPU5GqkA1u0BXSmMsnvpBQdUULRO8qRxhJw8ugP0Qh2dOBbRBB2oh
o29LHX5I+dMVx+3h6uTnZDz4y5DnPpjg9xb9yMyuBy1g2kFBSJ/gkv+dk6G0uK4r8x2l15xO6eRL
99emK9XQZ1vPFZOnyHRbFHcDblDSus2CwxDxYEXs817rGKVg8c0ncDsC6PMjKVtpCaaj/xcf4NN0
tZudFAHF2A5IOoRLK6MVgKI9ecMyDr9dgfgX4w5NF8eta9EkSW1l0kkabBehsxvG0JUxKe4BPW+q
tETlZ7p4kcYHP7gmrHwFHJuEkxmc7ezdCYcSEHriqn6AQA7ljRtsHEEqUNETU8766STG2W865uhx
BeSoZbMLD2EV9nzMgREGDTK886IpKL3XVYkHOPQNNUu2xNFQPI7rN7NcfK87SXN9txxKOqN4zUpe
rsbS5MjyeLYO7MHh/XnWBbSiIxEEZfb3EZkj3hRxLmftXwOfk86mFfHIFfZN0yMIuOUYouk4X0lY
JKRj8k1qXeHjbHCpPPTo03ZV3UXJxKwQESOs/lZaofxTOxpTES7OV/2wqv/aKkyQJ+TtBRmuXJtH
z7F55jkNRZGf+fssx8eyoAHZaxkLO3EkJmFffjGWhbNWyFDl0iz45i7x2dPzJp+53otO8Me9jwVR
kyej93OyKevBI82itsvKPoik/UBKOBcOCGQ3jNZVNiBiEaWIROXcaZV5C16yy816EK0dRhaLa6nf
F1bsWkihY9ubcuJV8snUabUKJSushv8+IfXsKyDol7snuznVJ405ChKqwhMJLIZkpW6tgYNx3B57
EaETFsToknAO021TkcX96bnZgm9EG3zhUammXtJIxFQc4y/P8XeUwn9gGBhKJR3E4wjefkD4e6g5
N1f8mrRU/Zb2GLXbleOUIG/I5H7VJ9MXUZwyEGjG5YrDuV4nruz0nHhMC/+F7RjWYanyOSn3IjJC
MzUV819tOkFRze0Rsyvu9HP4HGlCt+RlXrcZFO7eddnNs8o2yWOvLNDOqdaCiWEKxGLMERQ2kuyD
1rU8ry+GBVXRQ+U605dpPl0FhER85oNvQxbPEvjcbYfJd7tX5s7ne5HnvUjgOIBNkitcwVF6avbI
sGHyW0ibk69+voPiJeNsu4Pih22c4urGs2BkDlK+cAJQZgDI7LUp5HCnY9H/dcfoAqnaDghFvu+t
ngjIHuniFrWwG82907cYmvNxhikZe/plNzeslCWzfJaHrl44DSmNcbDPFNuJdZYjWDUoVes2Z0vO
CnAHzo7ZsF0XiGjUWLXUAEbQIIqUt3FZw2gf//g1eY0WVGCKDQprrvf4e1Dl39StN0Wa98tgN2h1
NfTtQjnmYDgpIyV7OF6rO4xN+1TK81EPAPjd8Gl641VvL5gM3s2XQlm30tOct5Lnk4kczgTXeQl0
axmHVroWkWNblLbI9ezgiGegPE/1KJEhsj8EG7UFil0ylfnurCE6gvhA93Tf3zxizCDlYXY93Ozb
Dpar4bpBV5Yf3jOUdfcwZEC2TJwW9rYRUZS9un7vK/lzYer3rULzGRsuqTJH5VB2z6q34LeQM00/
9PMtYUhsIzJrUbwEuzc/dbHCv2VGGGntUzckrkaKXa14PR7wdD27WkFadkU23452Ep+NlQenQQ+p
ou48C9H4UDlZB2c8N2rU6cAkhIEmJ/eMYeau+MpBkL/lRXuZDPl6+sYwvwJ9DrRgKuCMkzDo+XAj
goj4LNujKmbyiWvmVmC5uX/iBNbPPPvU5/6omqyR9sG9THK2mkFb/7Q1vH4WOOgp5RjCHfx+8an0
N2sAhLxLjyte/vmfZwHAbr+mFhmuqg/A9ML0C363Tg0V5Qym/1aURcTY4/+Up9m4ptNt6wuKozsT
fQXEKMh12ZSLkhJMfuBHacyRr8s0PyfYaTpQ7rigztDsNTBsWnSXFQkPznIwEijmwLzx86aq9iV/
AkykGKUY1cjvtie9e5hCgPlfMiYjETjGL2ec46YYZqS11TVZJxr9OtQRBE3GTb2IrWRyuZyS3gTD
5ql8epkO33x9/bCWtvXIzUejX6pM57yJC1CDpt4iCbiR1Q2jcZmWNmmFKqckm1YsAWdQCoJCYgEe
5CYIt2Ko1VuE11s+936zoIdWOy/jHLvFrWeoX7BIh+UcQ6oDxPCYBzguBFde0Khb4trDE73uMsse
YZsWthWN7U3wCfxCi/UgfHIDfEW0mIkNDFZCUmSR9B63VDLCkSnDvAJVLXMTnYymbJjBbO9wPWmp
0DNxyEQGNSoJIJ60/TaC9qvibv6Ewv707f6aWSALLcjrSTp8gAAP29A+2UoVhScZZjqhNFYz2sbx
ip+hWMtiGRObivR65JvQWES7zvfE2KT21MjfLljlNn61Nad13U0zvcDwM+tZIgNxMT8AwgY5zIL4
OBSed1tSc8o9OWsZXWrsux11wXMl5apCazYAMgVzonXTTXrDW9GyUTwN6uS8f6WneDLMTQ82bLX9
EFP78PVv0r2vVJYRuWFnev4VlnFkoeLsquVaEHZkEvToPpx3GG2N1ck1zp//fWzKXWNpIJuAZALI
zKFk95Z/QpfS+x17CYf8o039hOe1X7oXK2bBSRCs+vnjQRe0ElWTEuhYbDxmzRdYC6rReW1wCcZ2
RgeIEoZ9+wIuH+KcjxqBDRVsmgVxHYwNInSFKNHFgoEvs0G2/BlBsqWk3CrMJHk+yAJ0zhufP79e
jlJ4hOfcWGu2G3w902+PffgukahcOC8v69w5I/zict+zWMDU4Pd3jiwXfC6xHp3jLZkmlYij6JbU
Q1pcxsqd8/9dcHjiNUm2FOhTXVUfgzWP5MwFewRCyHQQ9LjAmHzP33rf8kXEg8l4XHUY/wELzobe
GV23fEAE+wMARFiTwIaBzsA8iYfwIRNQSRI8wVJ4pk42/X5cQg+rEWPEtUSCupEzsFPu55z9TWdi
NB7IxDpAimUbT5XJEe8CgUS9ErFCrZl2nYUBHYcAEJO41bPLBWcWBKjfajEAA2wxHYUy1+uCzxcq
RVBNCEI6Xp+YGVahIrU+dKHyi9+uPcBSa8SvGI8+dj5o1t6XQijz9jJCXXWBGWH/Fq6j+dupdvM7
OkJAM+AnzJXyLbf54fXvn0udie70SeLSMUrBdvkz30V5AtZLRZGtKzxKBz1gYysWUJ6TNUvGGcRY
Igfi1J4wauWlO4kDQ20cU6hL08jxTyosFaoYvnFUr1ATw9N33BjoldQLgUXE+PdvtBH8uZPRgdV/
Xy8r8HCz1/PKqULQZJEbJDtN428SYynKN0CNO24fS3df8iDP4omW0GVtRjsOwA/MtOspIgIfsVD1
VGa2eYEvSCcUDcv0WQhF856PRcwNjehxNgBumXaE3FdDAHfLLvS9JsCJF4htfgTsbWNC5AhGP38A
YNOedYpy7XpgxXeIPih9N1Te5xpIpvrOLslVsajFMxFsSsX0NAMbZYOiliqxMDoSfcKH0hf6HQwe
VL24Z+X3grpd7jIUWItneZuLV48FoyPQ7yvbkoDb8/XsHJ5jeUzXvuMIdg9J4gttMyMG/R98xXWl
gf48b9XpIFNYSnaN3zlpClUSde8WwOGN1vrlv31/PUzWxexZtMEQ6vPC8VIwOxSCLuZlXzOpHpUK
eHXbfkD2PHK/yVloH1x9Uq5tJydH7/xe0La9GP8cB/Ck/0RHPS7zuT9bldCCbPNxk639MMK8mrw3
R0uJcqnlidGCqcSjFjMHgNUGEWlzbFl50jp1UzheZaknVDmlM8Uypg1JT81X/vDkKjU2clnkb2+B
ZyBGu3Ofob7m3/PB7qxldVdc7TrTEbnlz+Jr5+GX/6am46yVwQTLVebD78W+ej4QfZ0NtdWTjTQ4
f6BcF3Ee7rzJbzJpHj0scYm2DvLCGNie8UxdItmp7VAK4nqk+HeIdKhPFZpiFsAzEgx5JAKH7i5M
+h4Wjvj3nKIKJfxXMIfI6pGxiJim9OPfQuedkiAGdfpsgphdXQWuKloJO4d1NhpYWKR9O+ePdXXM
JkSACkLz3N4u3sCAGTSVymbmDGZHR8OCqMTbc1jnsJlGHEHpTAc2UJmXDNnTT/RpU/YfbjoF9ype
ZKbfWiERlMO6MvYzZuLBcAH8BiC08elz8febnEiLHlgN1Iu49420URbN6zkI/Sqsi7Zxb8WXQ6TD
eZG10ZkENN2isakIU/xNySD6R5VkrQeZpIE1V+hSTcDyVEt36vQRBulmwasivkfVw7AEIetwyUpr
hIw9mPSHf0ogsNSZddWZG5+A5ot5i0s0UGKJqkqcbUAB2aoDfWiPlojEfB1b+mD/TAvvYFPOK4ps
XWst30XauQyca+TSaniEcw7MiTH1LKDw+9NdqiQzjCb41Jx+869IrZEquJ3p8CuA8fO1TEAl5yH/
H/iKvPyO++4qkZfSYifFJO+lwnpCPcnnGY4SlBSfO5W9xz3FCef7VAxfyHK2L2SxpOtNz8goKJiV
gF0405+ZdWdVcA34LPPN+6L6wVDLiR3dZvmW97bxFKa//SKzY6AoBLGvsQmGC6Gx7iFoYbJ8WwfR
mskVS/cn/hzQXClKSR1EZSJzX0DosIMuuuOV00KiAG7dL4dCHwtkabSISighyHrlKWpZ4HgWQ2Qo
7UScNkYwWaA+PJeB4qjcRtbxeE9v1WC9IiyHVjH9YBxINODQSIBoiTRUdkcSJxbAkGQkEK2G+KBX
5uBRGH28+dOXTMAU++i6RbIrAKkV0eDqLSOBoyNiSjvY5QMeryMNSSqbaVU4nygqMZpmsxy8+nXe
cQgnf1trpaOTClOp2yjgQ7wTsxJxW8W79+8EusaFBAR5lhdZ7EtcVMPF+E2LEvCc5/DmZlALPFxZ
y8W2m1yHNXfC8xPxU5RtwX/5U/Jy3n3NgNDUkhIo1MovLNXlNd6x84Jdp+uNd6qXRPMTj86Ay/Bz
iKYSdcOXAaLdivnmNRFBaODw+umKt8Jzf8F8sYo763ue6FCJIUFkC1HklVSwxetsm432Yv5dmDoD
wfeFpQln6O7SFbeYYqjYTSeSJv89YxPQJl6RA9gJ4s7jch9rM9StrIu5VeZeX/s8BYm8EXSUkHfy
2w4rPw9+Dsuu7parovhQvznny5ZjsHhL0SOJPuZ6RovMXqyUBk++f8axYb51sSl/66mnoxrMO6Uj
ihloYAvbe5LdedK8tThXfh8L+XYi3mIu6iMY4JfEZYspDFYBusDO6RcpO0PgOY3ngYsv0y5veVmZ
LSVxZvnItLZxY1KUU+P1Bau7bydGRKXGtK3pglabkhGHaSFaj3BL9h2J1in1TRCiubTxa6boiYq1
QduTITKK68YsGcgWINmiz1QmT3AAUCK1XDSAgU2Mby8D9eWncM/PJkua+D6iigEeSXqpRxP/zeNS
VYcr4XK5HugRful/n1O9Fk/gQxRgqbuTFzdWjPH3kM12vVRs0cmdmHl75m9BsPRLd/IaC8XLcKOq
al5ZlOd/MgwU5Js2b5GvEAN/rvczxoyvEZxCS2lZEiNJzKIhMNvshdEmRwnsVD2U2qMR/DXfFhty
Reeujc4Uu0rzC8dTcq2EkqZdaNa39hBC1Jd14qHn2z748zCgg7Lo+IsgxKKJa9wVX7ysYucmMfYo
DDkMZy7s1NGOg8lTfR95DbiyjYU5OsDHv1UomalUy5KOJUeJOxLI5z7QCf/wnY/hWXFTiHafCsaQ
Adytx8ID3TecPk1cmNd9WsgiXoZ/RuvhwmBqr0E9IP72IMNbJp8TAxAftOu6UzH7BJ3GVsVhuFfH
D0s5pK9so9ntxoRJtgXX+3sZYTh6hPxKTZdTMmnNySPfqI7NTyeD7Tv1XEvDIdLAvJKwYdmK2sBe
pDGmx+p/WiJqtt5Ajwu3TnvG4KozHCT85FTrWkEEgWARNlPj1nf2weU0GBGPzyQSgXWCzoYTLkhN
tbQOdEVpOLNVDrjMD7kQ6kCbGxcRUM7ylcGVJjIlWlliso8fCEv/pTpzDJR++rHVGatXZ3Ahgcct
hXinb+33qTsRlDJDLfYY8u/Koqi29wCf4/uou8BtoRpcY8WEozFHQm5Tch4TrH0+YfwIqAD9bfAi
JCQxXOxwrhGr+OOo52zuyn2/9sHNCY0AOD6pMT7Unk8Z53eTZOX4wEqePrGowFtZd2Z14AgFk40Y
l66JQAhNIXc6OKfDMKXOJGx+jzv/fJaywf+OujKabUJsesLgD2vqCK5+/JLrlAMwnkLPs7dMhW2F
CHUwPoht2p7ESa/TxDM6BAT8u5rJPdbJbtJzAD84jz4hlym+0KqpAsnlUnOdX4HE8Auueu4/qdHO
KjcmGNA9/cJV35JzTSg0IlYmn6d4crOw+j34oUF+qD7vP/gqeKBDPakMdvc9sbHpWWSq3mVlqFYq
KzpyE+3nNnzBCkFHhLoBNiATES4fbYBZ1jX0nH88lYlvnGDC1qUssDEoRCVwuwS26XqUtklivq3L
Ogb7g6dGjLU5rbfmDPQF3cf/A5ikcAPpwXj+nMxVRSyEThvAV5NSngsVCYZJ/mu6fDwn2m7fnI+v
RZfps2yA7hVsS5ggjIuphlP0gWRVaFSK/TrZn/hjy3I/oOlmZMKvM2yjM3LiZkTEH1lAx6O1MkxA
+Fwu7wARvXSRk2CU9ml8337AUgVHz3mTSW4YaxA598Mr1d1Fszkd5B7hQn1OvmOcG5jMqbhz6k7s
24/GFH0M0xoffT70ciItCIsxWy5+GasduL5Ggs3cpEo5mvlzc05s9UHW+YCaAF4cC2kasDmOGOQl
xhADQdiWXmpF3wHCcE5PuosWWdubemMYXZlNZ7QvKCWihn8kz8U/mS2b5Sg/7CisAYJ9Bb6WsoqU
kp5mWvyt5e870mHS+F8YL2bzW2SyKoe8MYNIZAA9fTLN7NQP8xQu0BXjAY34IfLsslmf+qezWjNr
XsPZdL9uWpRxweemhEyive/wivWAIvZyct6Xfe6xkBHquq/EqRdOFn0XI5HVxERj9XjjpNVe/CkI
92VphD5MsCnuAJJiWItBMgfH4qbkwWSWOh/Z1FZaZoqeaD2ktByxAl0PvNKDNR+fRthiGtF6xGZW
JAKq1CPAAt9BVacScSS1GpCUREm33Mtg7qja69XzEv8R1Jpvu8w7z/q1rK8y5Em3v+sUU5YLh9wF
Guex9T88OfVCh8NUL6MonW7p7GNPVPI0sQvG2uec0F9mF82Dro5ga1khgPCrKbqgmRwlxrug5lmg
5Y3UI9oBNFf/kojwpK/1nUNq4mUpiPE+SMbZ4CSmwKk/pwvHUhBugK9mVwB2ScxE3Igr/h9A4ER0
0bW+MMXAsZUY8yPTUnfZ1fj6A5cjm6vqp/8re1j4GcyWA/h7futmO81qvnoysJv54Icz/tzEdPGi
JsafWOOy0ah5zjrwfK4U5JgseuVBCuTeMTtidOTS3iq8EyWH18Y+vpI5nRaIGitYUHrTJkunVdqu
xLR2Am7gniAF2y/UDClq21I3t5Ff3EH5rRdP1zqarGS5TqwVf8FQcZ6KWhGswUUN564JnAGNiDXv
IiuOYuwbMWuud5UAfDgp20XyrgUZnY6ureXUTm5AqUECdkKt3U6rwY9q4pL04EqOD6zJIcFHUGPh
nl3Ei4iqr07pS29DOGDeFLmuGrzImuFn5P99/4H9tySmsX8W2VwFnOwcxo5qfxAC3qaaTCCymaLH
GujIU2RRQBX6ZBH4drm1av4bZaITnWEHZaaV1/OUyxXHyRy3JQnlQ7ARvCvrET6tBKd2Hx944O/5
oGsp/5B9t7oM9fTq+XJ2v5jKr3XmmyehioKwjIUey8hmGQLbkM96CFF/9YIhU+Hw105yvUVWbxkx
oLov+cXzHP5/3s27eOhXSMwqgLMyeUGjso4lu+cRMq/cEnCStuwNJuG/GfVLpXpsQow+Hl/a/Wd+
ppwb+HwCK38fZeuUXCn4FEVUZoLREef9TGbb/SXwUBxnGZPqzRt8vUJ8UtrYnG92RT5OSI80GlSv
+lPky3L37kFEIZYbXROH4jeYzJSDNGPFRoz2mc7m0G3fw1YQoE2oxCIvY5n7+Dxon7JP/y2L3AB0
fLo2feimr/8qcPZygE3jWw6d9rJTCj1qxhqbQf45A2MjhcNZH5fWpDh0exTcbr2099m2/SeG1OFs
YbRlBpjJnIdoJzgxa/oK7Vgv2p5Sy5EpjSk1fcwmwhq5MMMr30tKlaE/ZwkkIuFIYxL199xw+IWl
yTVtRCwTtahus8Nc8YUBFfs/l36siIvAjdKxbSssPgug8q/ojPBEdleYFqQKCSgThJd/L9WgV0vy
ScPz2Zv/xB3sB6J9Y5bnK2Eyyfq/U2yGS/rHX6nCr28QCAG+EQJ2DtenPgF0wE0Wts6hX3A+CxUR
H5jG5cq1YzngpDKdkKZH4azOkCdSfIQ7X/w540q9y7ehmNUnm3Oc4VX727v0yJecQP1IJP7OjQ+e
lJcnMcvB991nQa3J0z30HWubcyIby7L2alUTF4rWUqOg41mdzR3p09VTwR22xtq1jhHbiJxBata7
4qt1KlQqB5TMRHQHy2cPyRyHg+FBGpxtkWJTt1MPqfojMp0rD7pEwERGjcIdUX1/CX1mJMndLFyO
V3GNWwZdeSyavSjr4tnT5QwohZzSQkjuPyrWNi/OPqLU0FHAYkSb6aEogRvOCxiNDXsJm56H20VX
IWPQRpGyIuTyROd4z26jAVW60XqZgPfMquVpvhH/0VVo7KvXMONc9be6n+AxMTi3dCbsUV030fnv
HLEDNx9OESlDLuTRwhQGz/cNLlXz/himvP5P0Yrc7aVUdrbvH5jefPmuL4A34YbIAHnEe/UqHF+D
d391GluKPnfA4mOIKXdNbDBIolB2JX2ZQLAVGFiqatUWHjukhdaHruHabre+M+ZARk201W3/yfqE
91AMSC9BL9j7C52OlqR4wogcW7q0f92S0yQI7iuu7f4K/mP489NvSDOrPNZtT5YuwUigRFWxswlF
4/2Ap3XRjV1Ao5TiEq5NZnbJKKLpXNPMNKMltbuf0VCzxloXOgnwERFteL3Ugrctp1r2yReg8p1N
F9Bp7UsceKRBsX/ZwIzgFEwcQe/Ir2apjcWPwATc8uysbmd+LXplz2WFtJO18j9pjWzdS9ssepZl
1fBIsOAHdEV52KbhD0GHK2QDGlon4jBK1X9c53Abg+JUReSTgtI0QKptJc6MnHKNOFM+/9wLY3+6
V4c3Zq+H/viDZYFQ+vOHaEjUq4z/GhrW5w1F0WVikfpiyvEOARiqDnv3EhGmLehkJ+En/W53ot3z
5sL8WbICt3r8WO2TQn+Uh67doFhxC3pGfVhfOxjceH9ZhwrULXV0GkicZyJFxIeAg2O4sAQaPFtZ
Gyce1THYNNazPdQKGKeBynEcPG+s4YhDmKYEAQsxXFRomkO7c5JxX/bMjWoZEo2dXaV/avcItx4y
J8OdKau93wkQp1g8M6RReL9yOKkQAbKh2GdfI3j4Q7Lu2et+8UbdReYVuzQjbJXIhnHLfWTvJgws
ngW1m1uc2nEpbRefpBDXJ8bZLeqbCs/0UGdKa57YYOjMHzfWCgb+jsQ71kw9R0I1eCw3blWm9K3V
rdkbgqK9F/HUZstVTUQ4ki3TEL9SQW4RoctTZlUFcss70D8eQMfHdpn3TAL7ZrmNxi2J1LcrPMNn
qTgaOZgQ0U5YqRJYoKzuUwtLHUzdvp+p+IE25APpZMcrIqDHn/jI6uQ2S1ML92IsyXD7OFXYYZKs
I8cefoHsq116EplsGNiL4enn3D8f0LQ0kN8xA9rckYOD7RBH89knGW5mzEijHc0PIPYv1FHG4WZs
HTqxGU3aHYpj1yUyMnUIGia+Uhal3Jam4oDhz9KTsSw0B9MScj+0pToOlt4nGYSFiUf0GoVjbepk
w3t408R9fjJ9ILBh+0EFBltSFQijtE0o0+5r2bOfoYA6cTXDRZADm6jEa+JPfgKurO6TKMbZFcEm
/77xi8cGH/yWULU5Ebo9FP01nhOzfqw+zf3TCKFzQ7x54aq9LaliKQDCsxeZTU4dYAU8TdpffT8Y
OLiMyCkl2Dq6yt48MH0l27vfbwWHcVqkeMPFAujOPjvmmCACcMn1DvzRFaVN35nEytyJMo4Uyxn9
BcrkRJXwLT5G+oJD2GvsOqxb1YHmgH3A/6RvOaUkUFJN53XFb/31EtlW6aWa83ZgfzHjllWxqLrQ
MOtF+umo0m1iKM1QeeYB5OtGGspLQDm8hOixLpmOsgCnlMAnfiE3doJ+PHxOH9rGPTuWAPwVkwUY
Kp7lQlkoN3aKVrFhoQ3PoHxOEs92UwSrnlVdT70VO7QBTq6Gd7sEt18C1XfNaKXi3HaBRLir1NhT
T123c+jLAPI0IOaBoNRM8IshZcvgcI39KoJkNiAOXr7GOSlmHrmcduAO+Dpz9DxuSQe4vbr/Mtot
eabj0sO6zABO+dPTCS4tskGvXruV77lzZXmPUMLqcSpv0e1W9E5WRhATyv9hcwOSIiyo/bcNLspK
C09l+wbHKHe+gHtCehNOOceUcl06vOY0W28xL28GX/Nh5Me/FGHg2Vg4+wupDYzKpHcmpUAVgVyZ
rWDvW88tMgO3nq52jYNvpvE6aPZN3yCKtmefQAcEoCvvfy6u19Lwb7vfGmwK/ric9Q63kNRefslM
aPlJ1FeaLwUvWKa4HM/eHjeN/qvlSXEKcdiTJNaV3mADkvugKpQb3/mJgJ/MvHbiuTwzf/7t681f
llgaW47CjBd//ac3IgVEBDGlvwUVhju79kFTQY9ESKCZr6worr+hbztfASrx4ZnA2MMo9XB9L17j
lbSTFrqOvoFR5GuMxIw8iHdYnzE4ciHxyIJBxg5ACSG0WYIKRWcd0OQmeTYUnXh7QI2TYkTejV09
gWg7WKuMAktvwxcaeYbY0PMEZB/jdw1FBQJ4xG9cONZbnptmpH56GEPeGMCEcGv80yPGvJXxh4kJ
PapQv271edLHxAUrlHZCcItXNfBHTvBfKIFfXKH+v/tj4MCoOQ4P8QiP9pESkKSVpPKwSHht3Sre
g6h1+2b4Ju0iol3TSjBUOcRyXs6k2hvTuEZQ4iQNKb3dLzk1d7ojt02Q8UC22kkRQhIzn23YqfTO
+khD3lEmy+Oixf0pXSADFqhhZlTjdNlQSjTg7F6Pjhe/kNE/zFV0CX876saj5uFoVTUAzu0S58Xb
SqOHg91KlYjQxPpMC72IuThPfzSCTqnv07gfBh9bXKvhvODSOAjRGO/eWyuX/RX/jS9uO90ShbnX
RJDSe/zY6GM23IQHTsZ0UtcxN6BuoII7z3NkDP3SuJrPRtPXKlUzAI0I0ORC7Ssfmlqr/TIdKDhk
DvaFiyLC5ODimbijVtu0Qi1UNdpJudkzJFKZ7wcLQqT9gh1dLpdOF7O6yGN9RqfQ4v2YFmFq7lKL
hjTB2oUgCWVlA3XOpEynGGBQ/UyprCCzbatQgNyPlhORlle4ERWve/pwKbdAabZ6M5f6ifnlI+Tk
eimZR7n709ED8SeDgsVlbYYavEDihrpiB9UpMXfRSgHaFM7qkIvb8nUH0YFUahdXvtSzYEy/9ifO
Mfl/AIJPzoZ6T6KL7J2wXWfk/bKifN6Zc6hpUnKEAlekC3KgBrKV53etIQBlXf65gPoxQYWZmM6f
/C+mq1vopYCD2rqJDCnB3XGRl4/757vXAM7mPsNcOybqISgn8oO0aZlqzY/xWuPEaUp1ExRPKCjS
3g2Jg3YpUdiMRdvjwlDgyfhTF7tTUoTZ3Um9gcz/ENDh4BV3eoW37rWqgj/RBGK9KluhWSDgKv2K
qzqYBXQPy8z+AYVsZmrHl2CeREquKvaLNpvyvOQf4AIxs5DknjSlB6dkT1lnLZBf9m0jzJA+9rrS
h2ho8HwGm5qx9fdGAYGv8GubMe2Ki9AYnp+mD6VgbaTH8JDxwQd9Kq5lit7QdCX4yDi/73iVvJl1
ZbLwrxp1ic9Edz9/M7q5C/yOZ52Er1LQwdQb5GKpI4x2vr01nUkMFZGDFuewver2IokPg5kEC+GH
jSCR0k5sqOo6b0jr2E7O2Ih+3TRK0hwlX+gfWzgjoFYfsWvv0bZnF8rQQFpblgQulyPeZg6tX1k9
cEoVLpIT/wjyqXB+klVOKZ04vrM84N1KPJh1w2lBCU8sBbBBjlyUbnF1gJn4ZN4nE5O2PWK+pT3H
CwhWlmnIMUBWx4Hq5az0ulSbsu5XldSb7YGLqhrdQ1ySN7/Z1K07uNnTjmlqe2cKdlotP6sTYP/c
RLzjTPyuKN6sWIGW//VXq+i+MMPmfOmbSCSqy7b/M+KPyUrTsHN3v2s/rnQ70/bvzhGZXOht9BRA
whF5b4ODcClHp2SwNqrafb7AKBqtshrAIacMR56l8iB6qQP1JjYOVEXNT1zAEyncr+mLqgii7Kvf
CJMhmWFlld1EpN7EwZTdKEfVCRPZPf0/mwwjpm35IFFPRK2txnCn9zxCNQzULYLMeU+HVzYe4S+4
+duf5eKiPnZjfeTegH+Qk0GrgdtEYF9VXm5IJBGMDCydlE08etxuGLxFiBZNf0FaiIqBn+v7lHXt
Jx8BlopJ7f8kow0K9eQyR0sU6ls2ZXlRVfRb9KfVI5SLQVr+phqNDzNrXhL+S4Ej7m83VA+Ye/+p
nfwuohTsJPJQhE/RwLrBEv2+W7bTqZKSVedOwOqW0mAnUMQYPSxQeRXykxF7tyDOS5cPzoeGkW+x
/GhqLD6kBTZ/jFUJwxW2yx+6Yf+L6LOazSq4Xn0CnHJKJVqVobqLhxE8Axm5D+fOA+m78n4VfpB1
w7gsgJ4nFtkefTrq/wS06+RqMvfjYMGNAO10kTCUXuCLW+SJFY9iHVC2Ge9iFFjjKkXs4eEsMkX9
P5ixX7lekFLLccMhaPag/VnchI8Ge54iTsYPs2wyrpassHsEdEt10G0/bMLNjz/+ND5mZD555qDf
GvuSHpLwsPuLviRIhxns+KhDTeFKcQtJDe8nnDAmrfx773Sgi8m7C420to82CobkvEVgE1zTOmoX
khxzJ0uKHm6Zkh/SwBRdKis/9Nv2uimrKzh+M2fXLPHUgt/dGSJeMcrJQOlHvLrgL5x2NxZVUUL2
ECUTHkmjg7Yw6URF+sVC31FJtWNBfgu00B6QV8fWUNrNEuPS1gPure2BRY+2/4rYSs8LUCHBwXAo
vmibeo94Qr9OF1llbQNwLQasQe5HUM1SOHX0vq9p5T7Wj05y5OFlyvkSpS9U5jkg5WStTcMDLpgK
rbvm/CHMNwAywv8eEf9h1Ukx1pPzBpBOBXRQjh/0OqQUc2oMdOJQliixnLqcuLb7odkB/Izi5RvX
LnOsfPGptZqj+D+8GJEn9+ISPB+4b8qFbw1cQAaqxKM6hwy7MTwSk4M/HtThFIm9Ko+uQUFJaRGq
cBMNEdzgh5JtU5G6INxBoKN4QoSfsfatdE5/A9mypizXc56bdXjJu9BnJKHwNQ+Xhs4els5z4sWt
9HLVB3b43S5rQxIoFbB9DmZVeLUx34iSwSW/OEkbjTiCYZUTWru6Y6AlMmlx20vS0WTrDVUS2KFv
bGvQy3FkAbV+fPLxBZiuPnGEpdAhnHsExe+dgUvisJRHG0fIGlYuqBodYeUNWuwmmcTACFxZv+6p
gnIqRPvVfvEt7voYYrVJEfg+W6MQfGLSVbIbfyoYRGTYPjSLdDRlQQM10WJZ7uouOMW3QpLDmaKG
XY+KVMMjyjsGJwQuawtRglM5089kFFogtQia978OEVXVmjycMh5JtCnB6ThEMd15FeX2tZBDq5Gr
koap5l7ZwStg05l92z6Mk4bCQi+doSIPBTTGJD9NrXk+7rYHMxI6w/+zabv+RjXtGXX5FgB/iSMJ
ISjER6e+BkijZ4O+D1Rus/4389deePThxXse1QI00CfMGdWjKFBK/+5QLFKbq5u5XGdX+eno2VNY
0ziqt1TTyUOJEOIrOw5eOj5QAhSCk6+97ndpmtXSxHyZyk38FlzlLY8xdKTyxE/a3DnOpQ0/Iqan
2xyoQqle5/3UFKempKuqlDhUg6erqcOZg1XxcDIM4ILyS24TPvsNQTt2MDyWeUdEdHp78e+DT8mD
k1dvZD+dzkjDQRdzdTyHOS7kZdXc/pHsRLwtDmuSTbTUp7oSuOzXgTnZbSb0JNmqvUKbau/UkT2U
bneHgjfQzvBf28HqHC+4BJU689AHpCjGx8BW2AbgPO+6YNZMXekOzugPSjTj1CSCj9/eMZlXUAqu
fPujtjhzAG8OCBqPH3k0jYhUquB8A3zRRycWqCEQAV8+fUfcbFfvNkdGIW6EEfjKwOc99JOIaOAP
LAwbwLqWGCJPpYV1bpU8fS/CVG/xWO+YrmaBnNhGorOJwPJMJy9AghIz9ovmpv+W2B9sE1S+ZABX
3Vbw3Gz+NyXAxeQZtEPRuF1dMKiJq6VEK9qjjhDgv7lHIs01tJyXKII/U2QaFSNor1cxKPpJfl/H
T5BlKoiIA5ZH/e0RgJE9KgB9hYe0mwlaBsbBMUnPj4pI7u8l43t3aByKNBQPPa9LpPVDLTeReAe7
kbrlMO6lH/d0t6tePfego/5trZNM1ca7MF24oVM61pqQQ6qI1asbwktKoaSrVuKJzejMvTZ9515n
jT4oNURPqdk/112840yCcrYHoPUIJT/yL+jFUTVyIQ170O1d82HjAKQhq1hkv5JwH3UOibiJUZJK
dr5uLLMlFHbG1YMT8U135TaJGNRS+TyUYAigogGK12jjgzpuVPNQCGy8vsZPtHYfcnvVYbs3B2CR
spZcjk4RT9pzdO1DaRmGZhotg/bFMu8kGGD/HcOpu2eaYYEiQPgsmj/IMLDStujt3OI8C2FZJMkj
xotTboVRhH+mI1KT9y6rHQwMahQczp5VctUbmRqXIr16JYDWfhFdiw9LmKAuCP8+H1LiXTkU+UTj
57h8t5iLvuxIkW6S2zwKunkysY5yrldgTa0ErkvVKPD0dBIDR0WvQTOn5ZPF8wbFeBvaCkk8mCW6
5TK5iVwHMVv4Mi6YkwtrN+xs8FBytRMtqroDWwAus0KZ6oSjOiBC6+OGzIaaN8fbSsLkiZxd7AGH
e4diWfQ+3a3x6I3vTKwv/FDQOT2iZZcm+A2hdhDWe9lLK74VcKEK2UPPZ5GqPMc6Fd5/8x81xY9e
WmwGvl0PyZDmZdr7FXCs8WyKbf27pVmB22ApDvGUxnpqTVinR/4mzRc7tWaECeejeMRvSfPZqJC/
mFu9k1yMcxevg/XczHTW4JZZmHPV62KnNEItpAdyRr8xw/aLz2lzflUVzsUjCsElwCtS1ZwXWHa1
VkEf/SOul3AZ5/+7peWUbgC43FwICcNtQWAPCM0RztSN+R0AsAn2PEbqnkMt8UJK7t5cc+lrneq2
+52lgMo1V5WDT8sgbIDYwiuJIPLHXy6ziBqp1m6f12uYF8EOpbVzML2cYZd2zpG9kVWEOGSRSOB+
wHVu7Sul7WGr2f+VgHvusYioP0py5pCPwKTOMEvnyDk9eXCGlKr+lQj/2c6xJ8e29vJZCjS948LM
7kB8Si8fpcgWLQnKv9Zq5WR5yVz5sHhNpn9Q9tEY65AwiUlr92TQ76A3LpfmsS7OxyzGtluZqTNH
tUGet34upty4SGapwb9OTGj4nygMFFQtUcs95d8NrKHjUlxksWTBeUfw31uRrLR+xB9d81WD/2bu
2fKh//DRqmnIqSvToDpyXL3oL5iTcOXHS21SzptZmtWDwuUJe3nUnA31TAFsWKuI/apsnB2HhY1M
XXanBylrtlYu2kmRXiPXU19HM3bMXMcTMQ5wQZxSrBTiQLnoRNPO8MJmAPs673neCFKGyOF6pT8G
5SD7QKAFFvodupeqcceH7r5a51dG37S9SfBQAvzLyi/fXQf1PIGWDzFtOhx/JPFNuwpy0HRrH+9S
ruiKM7nNcLX933qw+tjimjIirEmwQaqznZgik1UT7g+3TV23aQKwf8yn30/ojv1g5Yq7nTuJ714u
EuwG1fU4mZSSnJAd6miR/2ItqUJUYJNfPpPXrbbVLyQ60sR8GDGaGnVKf09mlbw/NJ/DHj03MM/k
WB8JJAAOuVI2UmIE6FMnQS0Ksxk4xvbROJRS71gXQqPpOPO157zhGxPDXf4TyBuyLU6xhMMw0KIy
iYu9QHeICOL0CeBB0c4D0n2LdvPlXUQ90/mHUOqP3HfyYY3CLFyxLRHbSzE361fFk/B/9EEqZcMK
HqqN8chQEyP+A5B2VnfXsJl2sdjFj1jw3QfD9CsuGoXj9LjNidpsV7X6eDJYO8q7fspbFAI4GQTu
8gq+5eIRsR3jjbbiowNqlCx/UIV6HBsris785UKnbrC4M/BUfesbC8TagqzRvvaAyoxQd5mQJBcL
OvRbaYhfKG836WT8H3dZ+fCqZJZvkTIjnm0yVjorm2jGeTNX9eamsCfpTjBLalxyCRyKE7dwfHba
Kik+e9+NLs4lUgNs6npn/o6MOZt4WGrMP0SzzUKyYLa/Wjxi9a25ivXkvaaVnot3KABZT25JyXCG
aH7FCxEPpQbgpAey1uz5KtjxJWrkuwDiY9ALQmOU5u/RQlWMew3bR6XRTWaCSXw/lN4s6yi9QK+3
JXe/ANU49/WemtBdd5wE+A3G8+Cb934DW2+bLyOBR75L/Pm4coweHMC7M6wt0lyHKX/F/t861YOQ
6pxRM9Opi/ZE/ygRPtYOkeDDGUJIkC9aklQnmLUU2cVcoPjwguPIY7qvZwolhHZMc6OzZzYDHs4c
Q6xxIqYbu3lFK2LDa7axtvqICP9W81EOQrZre7eb20VPx/sRE6oyESinz6b1gVo1yAgxYEUhi6JK
IUxFte5POuCB6JuE7DIGh236aFExcHqZ0249Uervq2m1FG0aGBq9A7KbUiFwUSzY1OUdabAtEJl5
LxFXX/2JWj+oFzdAYWZc162uC/fcpgPyb7rzQ3XngDOK00IwYBJClGOvrWfodbh6brXqIjk6xW9Q
Beh7wyoARHofyurG4kjvRAOdXm9LLba9iLOTYc2TCI4RLKadLNe8d7W3Cy4bYQVwIa/5ElHq3kNG
WCUh36CShXdCOQk4sJjnKyVhz+uYRpNl/vi4y++M3NRt9vwyC844kreR6O5r6J/syDULAwH8K3d7
2WTdzHtM7An7t2hZ1FIVQQVjRonjLYO9z60u/r5tGekhW09ka4suAkpBK5aDQUWcsG3BbfOp8QXP
T7Zk5aCXfT28vVY1cgcCsysvhi+5JA1oK9UFozMW2tz/uVKGvSRp2bagCwvUurFP7sF265JsstFk
cmSrEYPvXTqQ8VepMpefZS6LIOS/unjMoj3xfpCUVZWnIMh6sgSJwIKP84rWtKdxxWLtGcaH8SJT
GxnxCGaI+GZHtFfy8TzfJoANgrwLEF0kJ8OAL4Dc15AGHOUQA78OSna+8f3rwXREQ6phzNtoe656
T+nsNLVByF0c+a9YKuXdwtFLjXJLoco3K5XwWNHv24BLQpLil5vIh1qIAUEkK5KZWpA0qRxnL3Cy
4H+5zUuTxHZEVbE+pkQL5qmSsVm7oCgPZ3ScGxvoIp16JwXWaOZrYtjJEKghtrnouDgB4obcD4L9
xwYsp956QJlLYNlIq35TSM7vPnmN2NMhe/sywY6BLy0XfXYH0i91WXVg0S8J/bvuttr9EMr+RR6R
cNaZZuB4pP9PdFggns77q7WSY6qhBLY5b00C6MznchTckZT+8nCMEnd0cdo4wyz10DP0teHrRYpX
GdBLMDRyEjbJSCQBfT2ogx9oi6SFU7TPASvMOBeF+u9j/RtK4Jg322CQliewnrNxjpvaXJtLxJU+
t968UZR1JEdmw7e7Y031UQhPh5e7oqqELclnhrBDAEfC3KxubdJyNP8aNZVAVWgnxqsrTNHrsF6o
qgaAmrh/3nC8htzP4fYIQCOBBBtGFTj0169Kzdqb+RBa7YURgQLtzlQx5a/6fYsYcNOpB8i0cEpd
Di2jfPhJ084lDkeh/xKUWDNgtqmzcnNCxdI5u+DiQrqits6onq0yMLC6k7RjVOILQ0Ln1Zf8TVdr
y5VoXZrRtMfCOjNtvw5OB39zDmaE0QmuBedXy43M24C6WNsdIn0Ra4rlivKujt5TcbmdJu2yszzY
k9d8jnzdkdzbAVtNTz+7OQhnD28w1k+citd6oDbwhbB24Bx1Bhg07LMLoEnWXczSg588Bd2T9PYo
L4pVHwUIJh+Np2nw+zCJSU/sCAB0q3AB004p57s8zaFytDyOXUtFnm2V7ldRgygCHnp9rV1R5LTD
MnPjL3lgHd6afVT2KUEuWNuHIuDJT+dNrciQRcOEWyy2TKvm2eomXESOZVuY4TQM7bWzvZ/aXVM9
+W1y5uo8RPhjNTK0b/8FmUXT+v1WveS7ozYVLOM77arWZu7651RZXa7iaK8H264YJqLzNHH2NReA
5Z+IBAqKD/V/OFFfBYtuQNt5jnRrdD03a8dZe6BzgfOtzYJcMjqilFe9ga22WquE1lmqdCzuQ64K
ihxkyUpHi9KZbVne/i7ZzUMqQDay3WjpZ4vch11pwtp/ia3AkU3lZGV5yXRCjMWOSKl9Z48s1HTW
BJSkzbI8V15nm6LcFyQ8HNWLbja6++jrMuzOEtKbdUXTbv6QDO74zeVDmkwajR4G+fe379o7p44N
5gRhG0choZsvlfi86fv9a3MD45tzQDnmIS0RY6MQKyahyV8kGQZNX2GQ1Y0hmt0fIglCqdjV8XMD
p6rlyGZ+bFZUbWS+fWBe8t5KYlQ8OuECTlnjRa4UTnxG4SecTn3/O0wn0/j6W0TAX855jA79/KIR
xkwBI1EVI989LJslYuUDIraC9zbTPWnwAtAvT+t2mVJWe8OWp1KSCzWcS7odFK88JU4yEZf+njzW
PhW+kSSA+DC8KdPPgn0Y3/4p4VEIh0s1uwVC82PPkSjKb3F2n2oX3JqkQv42nEznUtofQ3PO+ugQ
PZO/rOaj+E+m5+XAu9tH2SIPq1vsFcEqQ0RcI9/vA8HjgdG8tzyqXShku30epFQtw7NM+bV+GTC+
ug3ZWdVppHybzonl1Mnsv5laquphn0zy/SnMCIpV8m/ZnBqw3LetfWwZksHasWvt5S4kis9wRgxX
CJWA18WsCjsJPaMVvae6pbTKnrVYxZ6TnVMG+/x3JTCWqHopXXDU8GS96TRqrwTNhXzz7Ul3Hcpf
pOA90qcupSQ1j+RTIOTyo3rwYctns8wpJl7H0ALDQplW3ljZc5SwaGGoY+SVfWlzvYf69yPbaA0i
Rh0scIHV0BbdPO4QUsNouOrG1n6oJJ23B0XrOsNDWSQIoEMw9x0DVftVKk3DtC11emZij3V7TYHX
9WTYvc1rIQeCBN/d73e282L8S2PQezHFHR0YTn1nn3jPxoNZE2kAg7P8RQcz+GM1c/jxSiTN5/cd
kGNghg3kFDbSerReSm5/tySUjiH5bR7O6277ntpIdVJthTlpqFj89YLJtMwtCAOHmSmF3hnE0MxP
jTkd471nC4gy92lte1zqQaqmqfihCCt3YK6VUTJb0K4Xm3Jp6uoKQ2ZXi01ne4MosimfeL3N9Mpl
5zhL2O+7USyu/6vx8hybLLmCqbk1Op2mr7zQV6l65EOsJV+WYeXbaWxnBtBGG4VH05dID3EtNgXR
b1NmZjdqEYAiHZOKaaOeY1sDr0yloSFs3KwdrQYD9MM/xEnxzgq35x8/9G5TCsT2e5i4hSlm4SaW
Vs0Jth7Qt3wocFeed7aPfGou5FHRhJpUxwTwnjQsPJnTvqarLYvgm+AlyofE/y9vbDBeHZ6ZjB6Y
ZuUDpI/t4QIBzX3iiQQY4fYDzQ12KuKGCdE/mUkcoTwlE0SV5OoTkk7pZDju5MlR8EVtZjNaYJa9
uw1E9i4yz6g4aVdOLH65Ff5lO5vK0Ziwar/QhjrfPAzIf5ObhMwmYymiglQhB8W23109LlasW+uk
gaW3/oPl8+ZGcCLn6MJY0PtkmDQKikiEKsddKgq8PNWUoatyMOg2ARn9RqNVKsTz6HKAYmJDD74i
TsxTzfhiNuE+/RjeReTgmedlKAKm7PtHcd1qlAFLjbJszm74P2F7eZmaTKnBi4ByXMNUwTj8hSAg
4eCz3YiJAkFsu10GCOW4KYSmCvAmV7yPignOHJBfLzNJ8E55HruxvdW7WTWCZju/tUBrZMOszyT7
WZMbEZuzjMODDDXmTLnhL/ceUuZV/ybzqDhEcmwHrpbgoYJ7hNmCTdQvvXXDwlWm2jk3QrD9qooh
Xnbpw9WnS3zz0kZvuNs5EkWO3WSUj4w2Z36SiPDFgtoRwf81r535IVIebndWPfJW3rYy3ZGvwAoM
iJmQ1Ikl3F5y4aQBzmWX4ZKUqhDO9bNRM/sb0JfCPcModDL9n6ssK+HEQzsFrgdRp40CoL5NvVoZ
4/0+Rx24ASxjUvThMTEiAbg0c3gRITf8JIVr3N0qRdzhYnZ7VpMMFWBiP4RPyS10LJQdv9Qie9Fk
VUOnauEvtSL/79LnBADQffK/KswBFJWaxeK0+sxc+Ojmmvx/WYtdsrsNv6izpNFBWEjlQ/InR1NR
6qrJdixFi4bUvJmz00BnzIfQxaT19kci85jMDaEfSyOC0BfJE/UgAa/CI67vGSIGAXXdGOTkFH/j
GTKEg2BzxK27ooyfovl6aZekLOOCBBp+/dQg9lSlJSFmZIpzSh8rSrGb+U0KQaIxNEwi5Cl6BzJv
1uVNK9cZ6oaDo3T9aPOE/qOgiUOEXRqvyk1FS3OBuk8pQkY/hAFNU2NWVsI08s/xn+N2VAlxA9br
fv0VaODai/EPkAWdsoKlrvONB/jJVY0sq8FfTDBjQNtRE1YyXy/wh/M6u1DddCXhuzg/Wfo6AXjo
7R2gKkJ2+vUhqPSWDETEvBh6GGE8Lk3lIBn4vYJ+QsYWSbq3GJn8lCh29UhEphsq5rFWJrSpodQ4
GdQF4aOnwbE07YW35wZausoXPLW01cLvfnhFxCvqe7cSzRuKCBhixm6dbLa/XUwIdOm4nlvBqftB
VCCWnYfE9b0b/Oc4BRZmxidVooK76KMzlRwuu/M/HgW5Is4L/rJcm8oan6ayz2QtodDI7clE80Xr
CmI8bNezdz+tNhOWpetos1enXuNX0OjfodXglNE7revJ9zTgWNBcPGCtGpwG9FnYf5/ueCfqpJAY
V2NinPFlkSX/m3PwLN2mKY79lE1YMPZo6lahWrFVBEqg+SAG5HjgO1Cy0oDXm9OjgyOFvu2VYiDE
wfHc2m6JYc58lsRq1rIZq8gP149d2WGLivE/Ee3nAnWoCCSpBXxjcFFZN42dZvSFHQK/iniRUui6
HR8o13DH+W++i5S+KcP8gFFAuzmMokcoCRP8JFd0DYpHYg51BcNohidglLXcdtvY4UzDmFM0Hvc6
rZwtizI8W7fmZrILC3weTDY8AkshUimyHeoBLFPXzflr1f872zSO1LJntWJ2Uss6KrZVxHNaK771
eN9DP2GQ5LjHN03nM2xIpOS82dQXuNcJ3KmMw5477gldGiVuoIVpSWw2N0KBSMiipI/WsU3kBj9a
0gizxTw1AamVjO0VuXfcAzfmlGTTgPQ+Id3piwywpqzk1j4BP52c3BasHY1rPQj/1XA6pN4icKRY
cTkbhfV106/Sn6L9hddnsj3z75Q+WEzCeonaYm2XYYxmYSxWn2cFRpZeXsSzLx8wRg6PMMkuXoRO
OtJVU1t1IwQQnQKEa3ky72/jkj8jza68CJSdWxKsTVeGm5Trt5WEZ/Mj7eRZM4OV8PX82v7MrG2U
L73/oYic8mxqREbWSbQ+Wtp2AFe/nvK6pcgk3GEf7BJsJJenyDkCBKF0F1aiTuMKA38jQfCtG3qU
qUkict427Btc4V7ksxeK1U5Pe4C3ZNiBh/C4PHMfAUZWYGc1LYjLva/bxJe+1fexPg+K5YPoHZsi
978nxWtZYrATTJBINWubYt2989ON6be5Bvhn0BrpJxPlbyoEcGZHfVK5hK9KjzctPDGrxfaKUYq2
eACAJUEMjMeD5N7bWHWylWdjAFBRyq2zSs2bhfyEWBHyq/XQ8vDw+sXfUUdHgamgZacvm9ehzyfW
RZd1ZFuXzGGP/g089EdhRcTzwn7ejTvB2ldnAHZM+YYgcd2o915taL5GWJTzWVVw/UQ9Wuh6MtB8
BOdW6Vy4uHEKdejTenKMqlGaBYbtM7lovl3BYNVg2MSAHpoMp8sGqA+B2EV5gnyDAB71cK5oPrgS
VrE2vgqV9tzONUPtUU98Mvm380/O7AIRpXOsupRHxcdedeQJVWhfoUxPGjC0lumRZcDat4AqMbnK
uC/d+TFvsPo9USDd18MQNZNqQZMIf9A1k5okVv6GfEtSMRNi3eqekE+xWtmw6c2rIcmEo4s9rvcI
UX54hBt0gNSYWQNU+qPrqzP+HluWC8C7k/Ys1kl649NLgGawXSPhb9WMj/Wmqbzv54pZTBLpqAD7
OjSlcarMngPt0acMMHII7L0ApTi0lHEb6iHFZE8tJsCbUyHqoHz2vtq2UTJL7QO5DktoOqaN5pCT
l+P2pMcgt6yTWQpu8BVfeB7Ocdbq07SL4cxm71Tu6TXlluvDnTDNArf6r60RoSAt+tzOBbAe7Nh2
XF0Gqeb6JJItQZxd3tnLRiUQMj3+B4wdOrAGmKCRRyabGbM4JyYvJ1uddQAJXFHK4WXYRN2U7Fs3
YzjuVFTF2Eg7xP8lMFWSf25s5cCI83ZNybYJKsOIgQhx5RE7iZn3JOgYxCEQ9345VKW79JCdhBdR
5/kDiv/gjdmTdQsgjlfZyB0B+NKRJ1KgRK3TSH6Dx0qsleRc7AP8JPyTqlat5V1RKaf1W4h2gotT
z8do3jMpOIvxkKTpuxl7Rvjhp02G03jTNO/Kd5hWOTwRyF5ujyVLJGVJYIVyikMnpO2RGbv5diuA
QNOvnJ1JwqBwSVVFIuTy16hqv6jPxwM5OjqIy3eIr+3+XvdxFr7xhL7OTYQgXXnoCuisXlbrjLfG
i+Yg1jbGrXpLQzVDHybU9E4ztmrZdRcEsQ1jtDSns7RLugis/DHJ5IQ67LPt8pG/2BWgLQXQI/vY
fVIFQp8Ra/8TiCFL8eA2rZV1pOvAv6c8U2VuWyDRBnRBFnOmUdNS1Trozxm7wQchOCOWk7KXEbmQ
CiuiLxybSIsf/GDIUcag9VNIxEQ8BDUswB8aqElaYYvKA8Nys7SOGdyYqcTjtxzuj2WEQtwXCvne
JKtELA3uzzq1U8ft1QX68x1D6zjeEz040VA5nW9w8M3tVssKF1fce5kdeDC/c1lqSRwqeFT+gMNL
lKpYuxDdxjg8s4um7cfk8Tk1t/Rw1sr4TxFhSpoFIJfoVguP6yRk/XkKLbyJFZBa/7U8mdlrrEqN
g/RWuza7fYmEu+pho5rFm/0dpqRgcmmm+ADZh0iDiN03+7tW4wbPXiB2gScsJsU+CBoR+TzORBsn
dyDneAZ6mZCsEgFgx2wnVGqoX6DQdI9D6Ki2iLQptbAq5ZKtPJ4fZzmjaCGLrCl8bhzwVr8K89h+
hHyM2pDZY2u9wi2hxf91ylskpA+oaekWXNXgQqfwTXSYJFWPyS/6t0YckjjUi6XKQGCwptPuu3mC
zfNOwOv6mgasFb0D+IJJuQUPAFIhjxoYpWOT7RpKPj3GrTiD1CS7ocIqsj0V+6G1dj5n+4pCVnZb
zDZPc2s49PVV9F6I92YgVjgEIe8pcRn73pCm8mX46NouVLmqQd8genb9Yo1e9x3TveEYnYP86dgw
TFALX1Saz3kvyGPTtown20Yk0BeCEZjlbJPYyjUbMObMxLvxg4Q/n2oUMcnSUkYmB/q36hMawyur
QTyQXm0/LjZSyTYM6KW3TpvegJ0XKb/m1AUrQSIR7XWrJ3Tbea8rIwk3DkbwNq/fwRgwwtY5eP3K
9H55R35FqwxV6/lpURLjiU0xQwKoNssyhpXDCc8VFaGGE5bIDGb5FTugc/9H6sqU3mRkqi6J6aRk
Sns61sAEDFLqORGsaKfW4hgWtoiEb/q1cLDOhPOr91wyBI4y2AcrNIwTerC8bA3132PzetCuAjq9
9dki03pEQK5b8Ohk5xkMN1f9L4cAQR58bui94RYG65wUykMgSEyEYKWuhT/WJhkCQriuLQuzY6XE
ZdMZULOz736ChiYBg1uDdm2my77hXiCf/xjgnoQGi7ubNyXZQlxlOxJatlhpOhu86o/H8uAzUENh
5EF+fq/I6yp90L+J2mTq+iWg4skOU5web7Vga1/sXosJFrhsQrBPR7YGOKf+zErSoWLSu9TlQ+Dk
j7oN0SN5XziCrapkwIdoqs0x4w8oEbjyilzny5bj+CmdyfTFTbjZH7GJt5JnL7punfKnGuu6L2vF
kTaCP2LsgJ0MlZAmKh1opVkBU2hQXt2lJnnnkdNfcwG1GPf6BrFXQQf3ih/YRNC/NYnFGQxhlH3t
ikoNyVARVuPqRMOiJ4f1yraHsVSHhYAm/whRIFfTo5gDWMSPSD2FffV4Cw3Z/Mv84wP9h/hDMzke
RGvVNkZKQ/722bOWMQjf0zY7ldFM59SQrtz6/o97AMGFJYHGpAVI+Hx+rPP0HF6VL99kecdOB9IJ
639hvpiUjWlaf79eJ1zXa0RQHNYZL1CKJmBqbOEjcUlX9TFzLAMF0Y2kUTU+5PWJm3y+a4d7uYmU
fBpy8kaz3Sgxr+ko8hSmOBOicXZtLKtYlOdoIy1yTsMLtOHgFNZpe3s21OWpT+91xbG0RC9Pah67
7n5NX4U7RBuHYYIZMsYmyb9j84KFYPp94DW6yCvLMXZqRiz3CBsNjhW6O6ktZ8RH1yzzJBbN9+0/
yarYDkyRuVTGhUGF+dVEmXwcgHCAZ5s0PfN/XTYVeqiQYm+1sN4ic8h3VQlDljfn8Uo3bp+OCIeW
ChV1HaLsilM0bVS9fF/eGxZpoD5f0vyNyUouoNuKtazfGR+OjQ888Ycj1oZXNbaFDMBwkoPeIlXP
t3xmvOJUH1iUaEpyRoCyBkHi6eNdj9YtWPp6XA9Qu+zEg52oqqH2an03yy+4ZPh4Y3RD+CHK5n69
diXJnVTrhRhLsYqKT7knLK+cxkU8Xf1iy4yLqWqnNCTdUg2Yh1gS/49Zm2Dt2e/6Eom8e7WIz6NH
hKKI5bPUKLqSrqXiTXbuREoWFcaNyw5A5fVEoGyZihw9+4C5rY1Vs1ekkC7nGAR/Q3fZhlr1d5Vs
Py2c0H54fpFHuLGrEumuoYbQEMw04o3Hq7z9EsJ/Zav5uR+3tFy5qIo7oPMne+23avj/DMpje+av
e4NcV35l3B3gdFbK5nCzXg7rBjMSdK4u+/9iRJcHzNB6Et/61cqF9g8QHQaGaV8m2LFYxee4/wJr
EnIN9eGOtfOWa0mwVYZZDHADglxGovg59/rbAnAbVZt9cXEm1QU2KcJdWaKIeboxnb/dgmrh7p7k
DpDPDT43fYeDZ3tdB2cYd2yLAj6OHBDs1+cXn//ycXtIxbQ2kx6v7qkbn5DruvGeeDIX6ozEjeku
o4vULtPbkpqNsBfGFdPn2hor948lxXxuRDMoz1oWpH4sqFGwCsnMOKbmcEPl0YVcp21zW/F3BrBe
/QQHXmzn/ppOkOEtKflFvy08VbLQK9o3g6WyDu5+6mE/D6WcRfJs4Y2FqxdtdpmjYWJMiBiI/Ui5
KUyoNtp7jVbKHVjuSwgeQYmNK6uUoldTjDqTiW/IiYz+cBMf8cNNHssto0PAW8r4teC9+aUQpVKR
88KI0hVhoSQwaajjPuHeUY5eYRYTNIYf9bc1Mkc5tBfBanKwlNo+rAmFHsTSaxcpo80ts7rNjCRz
izIEDjMq6vLPu3r6ef4cE7mtTsp8Au1R7xFLaJi9oAWjNHgN45LsAJjT44wA3+uhidwAq9Xh4Qcz
XDbHyfhsVKbjf4W69+yMHmqOSYKWJQdFZMyqmj1DpzR00hV2er8/pZE5ixP+9rPsiljj/mReUMXj
uygFzoCmce06yWj6rpRhVQMaVShXoudYj/brAW9Slte4ocqVq+kP6NZ0nqGrnQubGgLemxlRhyCL
voF/D2WLnxydj3bq00quBCY0XyzpsRHT6LNG01U1PdzQYsW4BH9LNQZsa3Q3YVh9yIAQ9FyqJfIz
5gOM09Rv/5HL0TCkZ4HJ3aGhIbKDXCrFwZcvjn/WukpqisILcbkAGYmdnEZrlxFlH3toWrAf0LU/
hPY1nhL9reDbLvpdfE05cocSaZeZfOoisN3rHoFdZBjIlqwqtUPDsT092mC4OJhL0XHAIpC9zXwx
i5krCaicrDQnz5/dW3Z4f+Cuscux+iL0V8Rgs2l84bGtS3BeOJ/Tj4uRHm/TaszzD2frOy6hTGMq
Sf7wYG54YNV6cda/xVXWK0FmRwMZfIZfqB/W2M68rSfS12SfX8mBL0kzAFR/gcVKUolCbsx3Pj5r
mBr0x4xo3N+5WO8NXpfcInF5QgqPnfVLzpJS+YE1SAXO0/DYILICoGjKzHhikG7Ckoe/YNro14N5
fWO50S8FnFLtgMoLQ79IwlUE+fgXwBeKXQkYG0PGJqJgBh3bMpjadY6mf+02XKB2TF9EuXm8P9sc
FSW+vtydHI9wQZWXs3SICsWUCw7QkaJQ8SL8HgY0WzIVsaDRjqCXHQl7JDlL12O6PCi+UAwlEvHP
N1/tKDxKRSxQSaR7fgcOLEKPSpB2doakDVHlUq1egmT1tYOFCoZQVtp1i96wqV7P37iF0mybKSPa
51jMlR/6aSJwSSv4WPYU1H6jsX1bD7gszlcX+asQxZcrv9O7j/QlZRW9PJiMTSwoln76sWydGnW5
gJb2HfMjqMfukEHl2+mI0PEwVotvTKmnPHP6/2ZfhSgYEgPIPO+3+6m02HWXwvIegABRsU0movSh
kzQJAydmqj51gcVW5i/fLeoY3zJ2mdMSm4C2zpKQYDTEbklNbAC4xXp0R6Ebwace5jfcd/lsegow
n0p3WEYcJwMHF8sX/ldgjx9ESkYor4RZIftoWlS0aHU1UfflmaBnIvBBMpMX4lcdq6B7x3Cu4w95
x+bYHxWetQnciQWrI+N4y2A9HJnSNOd5huN8T1vws4FVOkN7i2yds1w8ViWlR4LplaZH85Zvh7i9
hs2GyKYq2WjHF/77YPLM/Re01uZzXicJyatiN56PQux0JAh+GW2jLP5l1zDKbpOS7LGwqSsM2a1l
Hn3jEMyJUNpSaBiQbK0XoEX4IWN6NLT929wHOZLKVR2kJOWFsKjhDmFpFWWy34LBwgiIAgUZL7rP
T+id3s/l9ywG38ZamenCtQGIR1xiQ0Ktda6ArKWTYTt73Db6zY9oz5xDLLCrmqw9W31kjBtwpplv
cx7I7461KAfEElMpND29EuvUbFqRHb4we0yGI4SYv7N7lDfSfcDkL6VXhy9vlyDoKz+qa4elSQAv
npHm+2RiNaYU+a5KibkpB9RY81ubK6DrnvpK+UkuYyCeD9XGk0aZrSmvWaJkvG8UrqWLqjHUwCel
TGB0yLaXU+ohrCAZyrIuu1pPInnqj/aKYYtj2T0Nva15BuMGplctFC5SQOz56ghRptaTqsP/7MEW
B8YCXa5tddqloYTXV7ikftsPPpZuMln3sSf1OwCezhJgAJoDP6zZ+AMgVdNQVQFpbDNF0O6LEgtV
K8jDsWvD6a59nLR1mNt1uVKwsxcBqKRaAIPrxNpM6gpsCUAr+68YXHd5cCc4MvcuZp3+jVF1i0Pv
pAaCm9AWS+RqL7sgs8juIR45/M8Bce74S0yWO6x72XWR3Jj7WYX5vM4fncx9SyTyBhDnOasdE7JS
o9brYZ17ummhnG81z+k6QlK/Dv1lfsQ5FBQ/JBCAIAeU9pVnNmFWf2ai6jlw/ZK5awsd47LU4l0J
Wf6zAZ0D/YDRjn2Y+/iKrLbGPl3P0V1m554MndxWknQJCISwCtGu9FTmZeKN42k+7adlTwAy9clG
R10cQ7jgmpglk9cll6xi86BUOA2aIS//NX73PwjkEr5AnmAx7dROyBrCFFPvZsp7Eptc7KkmthYa
66icNOe4ApDFniGttgoOF6q5PtbkwIm0Q3ZerbjKelBkX7Yz1POk8DQFiiqpv9kgNepUP/h3aBX9
eyEcMajuum+bRBkAJwjDWIB0nOIl5W8Fxfj/td5Xap97EStdy9dWqAnc+dpBTzlQt3nT8EJZY+ak
1DQnFqjqLTFsmyfB56sDwPxLa+RHeKLvFZQdKZN2NSzJsOTT0wcS7dGjP8CkOqsKE4Vll/ldJJ5U
QtMkr/QKCVGof3q66+MlAn0pQ9hjVllEpMMB3rJ7OyD+efigDmydc3ckDjjBgSBZquiTgIxZIcJ0
dpy2poHd6aAaCSjXGVMSClgipDKMFv+zHr2gOSkaNGPhCCTIpE+vL4iMgtu1a6gzWOu3vQqtmP2f
jmliqfKIKcJxqXz36aVanxu5podYSB2lyqFXDlPjeANqgAGY8ulYfFsZ7TV3nVfuYVrq6e9YZePb
M8BZ0cX7RNCtvcxJRkwOUKEmt29lsUVvlaVPuotCu8I0rpNSoc6lyXiq8LVigDjA6aZcdYowILzg
SMsSjGofVKp3HF1TChSs0h5az4b2q9D+e0etIVs8KrovlxA52VTNYZbYAi3hcP+iDTrYpFlf84Tp
IrS0ids/zi8iiDIbwEcubOlK2cyUHO1Ac7jaBYT2Xggf9Yg2OsQ9WCdJQz8VR4g5Lw7NlQdrXxS3
W7h3ePBnpwt4myWGAPfLlxOVzS1DdXlyzJ85T868n8QBpdPrX5zDGLB09lAum57aFLnejbRqddcJ
DmrC9DxGuZdLHUd8HdO+yYZIOVYhg040uf1sge+v8sR+sUUt09Kf4Rkt3gfJ5CDqKOmYAfCW5R40
YVBaLbVQpWZmH9hXToesMkQkQEe/5OlN+coMxt6V92tbAD6+2b/MAP564CJjbqBJn6aNJhb8X/RH
DYIiqC202/TO68dFLzor12nSoPbvhJ0Vt+Dggzza+EvJdwg+wwSDHUUiV0Yv80U2Yta40KpYuawL
dMy1rpHPE0WFe0VLgzAYkJznDRYE8qkL1iJTjcV2eREZys4Syw1ImO0CQkVyngiW5ve8eJYMbZGC
jXFs0QyQ4KVMuv/abmMEfWsyHpI4MouHvWR415zNIfPD74NQJCBapfwGRfQOeLirgme9ezuLKdFR
CcPB6qb+HheBTE2AOkagm3nHl0J1aF9UOVwy56yWzbn2Ef6wk3QjenRLStQucztLMP+IMLi44STK
+/LMQH98GRaLPrsRotMpYPfZACGbvumbSx4HCLea1/js3vD0D/0PEq4zmXXTfY/YfMaAvjONBDdn
mBK1JeVkni7Yuyv467V7BtDEpYSKIG5CN1uVDo1cjsZ+Le82bYX3h9izEmmQdcUiCx4TCCE+fpLN
mFx5sDok+eAGCxj/RRTOgT6NotCrPdrmP62jsOxUefo+m6hKfIZ3GbgyZnlfYJiAwSfDS6ENLwsr
9LyRGz8vWsJprJKg9mgCwiBtYS2bVVfRmhdSkw1SstkTm4QlIAzaGW+6mjQJhXvbN5iLz4y9WyWk
O5yaLJ8UrplqLfiSQ0O0gmHMGP34bHJldOOnVp/0bpOQx4kkwWg7I5gd8MKerG2PW+ypKikz8PVL
WHnknZMKjiLr7xvsbZdXQz2yU8MgMyA4CyvIz4XhX2J0nbsXMvXzxqRxGWPGijDqJZ67Q5CJEOXY
mX270Z+fdxS792yOhIH0RpnR1nosuas0cWAw0iGt4RSmFBvyaDQsFLMbNFNy7E3KnnwBW9F8oEwd
GAQld+mPVSvarqCDXMWC9Hv47z0h0aones5UzMIcJdMMJl27QX8lYtWX37aZroO4RTuKJoOs8Gw8
oY5GL3ReuqinraYAM4nPJRARMsKkX2+B20HOb4ApM47ZyG75p9zgxyihnlQzKddpZGALKXiuJmdg
pyPmERooVIwCk95CFCvBN4m8kIXJMrMYU0IQf9FCRCZzZb2LyLM6rAJT2mh8LxMy/0nvbAdIVOAb
br86KZveZjOQ13h34KRNBw7UO4JJcTgzvaXwAJkdLE69L7rUF4H7xdsc+4k56+GdfiPw4AAqp2Qm
Qh9BJSCot8UK+ztESoRcnRJ9Jh4sGmSANGe2V+0GxmuvXXEDXDWG2C1NEAaMPS9Lt96OWGGoDBpT
Q+ynWgdvbQqQLV4SOCzIrBJ92YPdqpL8MwbPViapAzO6AEDF3I5BRXlVCNJGNRtEIX8SU9SGbuqJ
vI98iWq2ou6ZxaPjLJ7atvKjIcjHPBmIdwVQ6k66yv0aQWkv29Ddx2yKrhQ61dKGytoFo6PidSM+
/N82ucmOvfZHeBF5g8CHatPZh7e1UDbv2VEwwDiBzVNP4k4lBY9mAuB3fyYET3qJUQ3vAbVlEpoP
y0Nph4fDLHxPjmnQD35xexiRaUo2d/NsmAHWeQH1RY+INpLUS/yf5xX78896WXTZ6BeJnhvtFuqC
zEGXgigK+2Gy7XwtFBz2yJg+Thv+/1I4B41D2WUTziA6Y4CPDjbX3FF0xZH6LG3OKZNRP+7dTAtk
bXM/+9ipSx+bru+RdUk5s6kGoSiqxnXTknKE9zRRbeJxGiAPFtNDdCffNNG3gTFkQyZJYmyNg4Ew
fIAvWuhZJwzwJ9sqntdMQhRJAmco4F8FjDKkTeqNfpXGSj3eJdAHgp/vK74bk12qEFZkQ63PWsmC
puRN3IFOxx7HPLburx6sr9Zvv1K6qNAlFtAc1t1s4NPoXJJN+0i7gEyhaNqpG5bpX0jPIl2s0+Ua
+CMk/7yABgpUbMZLu3rVeAuS7QZbXVcKef9/6L0o4sN1KlkaQw4aIIpRKmJb79AvD1AYil4Mcv1Q
t0OCvxWPus2SLdEXbESiCDDGLwxuW3+OR8OtDFJaR7pf0L71tfk6LLTKWqVRNjCTMA/sVWfFZV8y
7ZZl/inPbRnvEhO+MXH5dn0c6TlxDYLmD6nkP3XcxqpOe9wr4Uw7pycfzEL2nw6gBhMki6BPZ1Lr
WDAWY+l+i0v4KsYBjEPB8SJD79HsROOegBXWlcztDCAYwcngBQF6BVflxubopnl2R0LLHT+xdaJD
pv+GO2UeKp77VMFWDVp4RnTab7uK16SZzcYlrOOSH+lHVbA9BMINcmGOMhbtmQRyPuj3P2R0EHab
95juBGtg1MMuvMrnYJS1MmXXlgo8/+TuRaGyFVjk6uIdRSJyyBB3DFZDjlZr5JH12CoqFcvHwvCQ
+0pR2C/wzXXUxNkkFWB6DGZT7D/pAjOaS9DsouMhI6jxBLFRJxajRQTo9K3qfbUONzg50/oLxjtr
KgS1Xk6GY8x5OgmDYeXAaXWBD5l0VjyJGvaYKsLzCRYJ/uaTmCmOvCypF262L9kA3eD9mqswJnPm
Y7Vj5wXVfVJjRxT4WVfHUu4zu+aFzn3k/p74EZxlPVVfLA3jBHRVaD1794d3nw8dIMr/PjVK8Gd6
ZZphnSiKrF7boPfVbHVRTB7piBeoIadtcAX3tyH8IdP96J5Sk9O2l06Ba6wrKsbWQk0eqbO/wdfx
LGiJxuwBxmugVI7S2Dh1f/tMdPHwahhFhIEk08eR85KkanqApCQQ1LemCVNgtUd/iuX3VCvijLS6
CjlHhkCrKWq5esDW8EjgjpSLAA/Pt4jrAmO2qVHwr8wKs/vqw5mUOs/QuEdeTN4AovJLu+XsNy0D
KBbPz2bSSRLDbHa1Mc0e/Dg4X2PZIenZIk3tRikNVdzNUU8Ea3Qp+t5tJfbqJP4dQO7pBozhSZrk
AHnIJ59VG9c5aZ8xqX1MDaLaGJUBN8r6BvXk3iDSEDV9fyUHV6M3YKdN3K50Se4pEF0x4PY3v5fL
hoBBoPKjMlfGXBjYRD4586ZySjJmaXSD6ZrZHk3Vtz+o4ZJICiauZCtgcqtN8/EilkM7wB8nH2uH
9vdpUyn/HZtwepA3v4bmPvqvRREFB0IZTWh80YccbGVUH1CRi20TEEGaBQrFh+lAKR0OASdx8krj
R2XKj+T96X8rq/X/NRz1zx+Rv2iHeBq8+C49shlGOAp4fHF+szA1G3DWg54Mx74HiEl3ii1TVwXN
VLlCsp5CMBjtdfNXiT6xTJXQzPg+UUr+jcNsijybGTKma0GFTI5bCxRbXNa1ItzQPQlgE9iUJ/Dp
r00mh1wej5GywVVgEfFKn0lEyyo/0NJgs5lRifUCZaQT79oFnxiuAbKrKKql37snUbg5r6qdqe1m
HPZTYm2voEaWOcec1VyMyiQJQ3bAn4OO63iEZcqa2wIIed8KaqJujfQVTwH9XAit1h7VhAde6ZpN
+E2brbNagjg6IfAEg5g0ACKYdFVsU49mkkUmt3tsGto0pFnjsvhtbg7X1f/2ThmhnCrmBeATt/xj
pqbBrOG9BJ45JhXlQF+wdCL3BPpkJlVsAzLCA/1Kyz9+PQlIQUepYs4WMeZ2h3WfukODJJVT8g6L
p6myLy5KmOucuPRF4R+53x4eieFUQmJVfiMpt+eCWhgzRYc56MfMYtwJDUZ5+JVp8cakVeV2MFmU
2sgCq1yLY+yILwfRijTSPY1RJNGOk7YsGRsaJq6Qxu7wH+pF/LZYbND47pJiDALbWx9GmdXqkN6q
XLyVZ9tn8cOgpw6DcGabLW/HEKKKlRsls8gc/RKknNX52dk2VCl/e8LI5cBM1qGCiQBGwz0AcAej
9f90eoVAxukOarQqwb8CYU4H4dIGyK7vbMyekIj+Ju5aVw1soAlSAMX7SD7i2nuUkgKRNjFg/lbU
qGscu0jO3a7MiEZtpx9FLO1FTKqsSIaQzqr1wXDA1Vn2IZmsSIIYscSz1BWp1soxeEP5gR+1Wg8K
iC5KBUL2LeLRW2y8gUmoP6dsAYCx47cRj8DVk2QcnP4Y5fSky/M64+ZcsVHEXeB9t95A2AuMmQNA
LTv1yoyAO3c1I1i+4+eK//XDkMypGTn8kudx5KTAt6z/5yhHZuafxmvP7ilJ9JeNm8p9QlCc0LlX
47CUF/hRnEpbSP2UpbI4BlBiifZF5MIJo4R2g9gJ0II7J6qy0fznfLU7WO2n0uuO8X8fXr5Rkm3k
HuKrVhEBbcR/8yny21kTDGmrKxnuMxy7zNLN8XK1NvCBIEDNNIG+WakZGtrwiXf0c854q95ar2/K
55zhjRSF+kckmwn3OBeB0Q65GETBPIE/jfwW3s0+NAQVUDzn7QbMaCOOwGjar8bzdlTazNzluOn5
2DTFkS00B6WP2HmLFP6jlqtqSU2PHZ3lZ6Wb3Hrm2/LBDLNT+haTThivXKRw5zWsWYBREs5x7Ik9
oxJdU4jR6tlU3RApPAronC09x9MIiwvgHdxyI1VEmZMN5jVbgHUeNQ9nICfIo6lv3TbvAWLopR1B
HM4W7YuRTQ2X5Uj9+W2yEDfoAd60o4dMbC5PArpq1hTCb0+DQgIrBvjtXo/Wt2Vxil4C+KRWFRAM
pvFmvf03DKKSz4Sg99UTdZdLE7LIhN4sjlhnhRYnHu55LjlPZSd461KQC1sACplnKbx3XCGXZag2
tOxhvqhF9xs3xYR+myKIvqcb6eJi3oK6DxvRUFq19vlRNXHtk+vRgX5RYzJ2T5OjYNnKndJ13gpP
nQLSPhi8NzgV4e8eTr6+OPjeb71Brbal14JGMJea8kY3TNkN3GjGpY1uwDCHgxiGf2/8e5x5uws2
6ZHubDAReLCaZ5Tq1nUbNE3CkGCD3uF6G/XGdZhhHKXkZSS/PFWge/Ktw35EEMSp3n/GDerymUtR
RP0/SN09e8mIN3zy1yEa4TkmB/2FaLVx0blj72Re4JvaF4oxnANCmGehagGOzu9QjxKRjSOxjS7u
OI1ppWSKxPoPnOU8hNAa2gk3KJcG4U8Osm3/+8kSZVBImO/vinXKHVdACTySprZi6tUradMsRszg
iGvwGOctpcvXlKUG+z8pHT1wldUZCtblAynKCwyp/r4VnmkKG+J3bwVmjUVzOkwh5Ign/V2uDzAl
xHUOT3aHRkFhV8uGjtzs5DOUP5jwpX9jzCb/JVC48E0joQchneb0s93qrop6vSLf9tGKP7VKgkYC
FYusLfeuB14lP6bOhtK+8B+bmnAyqVe3y+kOF/bnGYu78iDL+y4zYpZVwXo+iND4xQxb2d8B1vhH
VJJQz3vAmBDbcZofavHpBRMt9XgoFn7x1gTsNsUeP5gS09iCgS9+iP42Z//d+CZi5jkbt++VpUO9
QAhrb0PbPgcRXzHGizdLpP1yXGVINOMPio8GS8zt/sn5sV6cc04SB6vE9sGagesnT5u4avNYIei5
UqBQlIrAWaGXGbja71lUW87+LCw6UftmYRbuJf5Afn2HjP4o/woDorvVbfkIpzXmRwnRbjN0OjeG
XAsiUmy6BcLeZWDDau60YeiyBXh02syotieyMwNLksIu1ZIKcyUIbkuu31QQAhTYHr+IqRJsaYXB
Ef74eGCx1Tww5PBYF4AMqj84JcdmY9N8gMANIbeCLSzbTbYFS+DIf4ropggXscO3kBaGJm1bXxrB
rzg6eTEqJhI5gr+5eG2wwGNO0VWdIRcQSruXbQiEG6r1QkdtQoi9EVD4ZsceOTQI3Rd7JVnzw2/B
UU51RIWyXlzx2MsQf1gDgaV3BZVgQykGb9fiudjc/oOuVno77RbVjgtocQmWst3xAgThH/cBU1Af
ZBdgJ7sf5hKkOtjO214vsZ30ThQElfdsqP8uGUOaNh2MJZ1BFjxYMyUXbEsXPKHgAKjLaOlqnoTh
VCLOZbq93mRX7xoqi1eLBJPxSBEgdBzmR+hVE5JQ5T7cJQnvcIb8nI9LewhTiTHbVW2cKAedpG2F
x8UZzxWUx904/mj8s5MNVZp9CirevqCEvetlvm6tZIyY/yqHIZvZdPPRX5Xrb0SUVVUSzxwIF6tj
hK9fBHze/NWe4Z7It3MwJPonXZ9nmsDBM+ZYjkYRvkFXAM2dpcWJrD+PqCqADF0yUnjWOOdDPi1b
YXCjLeOtLap4CChXjFHw5dwJIGoqXtskJliiTWZWe+JXdxn5ixZX3SIIcwQcHl2sGim8Nt2HrgFo
C87dAZZXRZqf7pLYdUaoOWI+Fn3++xervJKbjXfRE28CdmYDzQ4+Z+HXuoUCuXebOlysSN9UL3qd
ZzZ8KkV6w0gdrMIS/m8mP+v5RtmUFei6GFHjHRSih6gVu3wKYRtkpEbKLOBHFp8LP9qdF9Fd91bm
ol6x9YfZTgxK1HFQ+TaXKnYQY3MoNLi6j7cG0TPB0Fcvm46kwppYJycZu0/qtHlt1GaiF8gXrVnh
e5+2Fu4Fu+wYSCUGBFLAcY05KhPPBGuOIFNb2wTDFNwExT2Hfq7Ou22og/8uDMyEGzsLP+ctTRsq
t3c/wOYj1zksR48TBzCiyUOD31e6SdTpMEvJdNJ34mJSfRgZff+kZf1qjJTLsBlDcuw6hFAl/OL+
89aj3CTAbj3cHicM5pNeWFmDBfB3n7U8cLoEXQzuE+CHktWw2RS+tfZTDL0HJjx//bUFDiTYow1+
NczKiUGuXAZ3d9F4y3tb6XKci8rUVHrIuCQiaIzr1Odimc7j1wO/7gobRWD5ihR6pHOBnubXmIqV
7pR4ytd6wmjP4O18M4dRM7J+8FnJcGrXTaT6uH2wXQVgO4c255AvBhN8Na9oi62uqVNx0FvoJt2O
P8MiE4jeH6XaTaQsYeciJd+1Okgd/JSsTA3gkWswB3rQzEZZPPmhtWr/1XNNt8VqEgt+2YPwh5Kv
J5EWgy21EPaFti4mOgld/4rdzeOGQrUUhrKV8erENEX209gM9NaqSPRtzMuIVjWTAwysz97gnsjb
Hf7zudzhhKM4V/dH1t6v3EJZpQQ40nUWuRRAHrvVqxduIN5DzikqYQSAq0jGnIwbJ4pp8SCTUDbg
qvyW/yuu6eGbO8/5tt8PX+WMmSBi0DM6Q38CnFQijUHo3nDwC1DHk8II2pK7zdW5UJSiD4FHVSjv
ta4LMiz76VOdnEIdBgfOIq4s2T0O7MjxAShWm1Xgza+eoZ2m5F015zwqO92bui6RsH5FlbjBV5wL
TP3qQ9tbVbRA9ieRshkuE86cddTorbHdgWqKPGZlXYRlmlOng6GLCk1zzsDIhzRZAJ+lNe9DA5H4
tbDRmJ9WqHIdl1r6TmUdQzCe5WPf5zbzluUH0yDv/qOwDmSpw9gsXPm07yFKDIweP4+ZJltMXk6R
crZ2ZM6B1IbqwlPF/q9c3WTFofFcuiVm9U9Q952joU11EcmvKaHZVDy0JiOfhQBmg9DJ1BW3vbc0
wVOvtOydD5iXrWIaYvu5Z+ikHYjYSVjYRdvyuouwQsqqyPgcGyDNv8lJ6aJR31B0P2NPFuwBbUwb
69LrSVBHcO+iD+euztl4B9bJBiSTkXrNnoOPQ8QnC8MQ7/zFCwt2d88CfJKh6a40YhiDvQspHWxw
J1CMGd/e4320azz1WgG4b4RFVKuK0QS9rJoJFU0bPNtrL+d2eaOLfFtu3EmrvytY41cvcfRFmfiW
dwhSsSX5ilSywTh2CplhEN0LqOCYYNdSpZrh3BHJ8bcrxzIVaKH+KdG/DFMmsIjbSN77ep7tQ1tq
DHvtAYWmTVDZOipA17EmJNNHpHjgbVdbTEvCE7J48XiEwe5O9Kg800jVFqOouu2HLC9DOrbfAmVf
Gwqgv6thXa7H5dAFfw1JGJylY/9tr2wBoik4yfafl7eXgQa/Q7ek5gFCS0ikKt5OSG24sSAHH/t2
KAX8Cnsp5mRQr70RmS5nFjcyVdIfe8IETj8pISWlfZOcfkZ5ILu2O8j716OmReo9ixNq18u0reE3
78dnQkoqCegd8yiSiVBpNIulnb/qppY1VfQRuQf73voIhmB5rWosM46MZQWqK2mz4JpZbhz8sgjb
ydBKZFq/cWOEBH7t96aduEpgY413DSQWVs3Bamgk++ymni/OzXYTZ92KOshZP8A8NCDJWKVLRUxm
+MD4rNxi2oxReAvEchUxZ4tW+mxy4eBXvX3BX0TsB1gbqCePrUIMBIVbWIzGSpIcT9ehRgIJotAb
c0Id2yIWBogABWvAXRpNG5YJ9+ZD8fuPXDKptRzg0a4PcEwJiTkjg34GYuR7oR+N9ZvnlMR/n4ld
GFPBM8F72UsPD2eCg9CqU1FsoJyPn2Mxd7rKbR2mu1X9Mo9gZQqQntEEkGIflfS+XFhV9iAvt0JJ
H9ovPizKhLOGchbv1xQFE5xEqiw2KEXr6y8F1I8UBi5O04Gr/zyHwwlU+lXd24P63KjxZrDI5HSB
HMhXkF5Tr5IiHoM7GRZbt1gra9CIicBT1albZP7trymbG8M+gMfDRlimNXjUg1T5OzXtqBtCfOqf
+XV43OVI8hXtRY10Zo+bnQQDCi1yUiimruSyEN4MK+csaMOXAse3vMD4ZY8Hh1yypETCq/V7Nk/9
FSrG3Dw8EjSl05eaRN9CFjeCgKcTQE6hOhCW4G3XpBBVxW/tkIKKXynBiijZ1O8hzlrOtEsE81Q7
TGYfh07+sUtTKS+BbndYwuW4R2c4D7VBQgGaVIMaOSNsQKVdxhJPGQVWON80tJliNbYgAQ+dD4IU
gVI/VyEnVFruBvbPAlee+nA1caRzlkLN3MkvjWQfO4qRM8uUTezB63UfX/dYFHWTUjCou3RWHRMF
KX5CjtvB0Ymp9kGPKx6I1wp2k6vgegLCRROPdHBC5qW0beMD7jTaBf0fybHQfDh2GYgZNY9HfKHf
f+7r3cuOFQU/Bwkpv2PRhTTqKbNniCw3BzvVCvcwsnR56hsM+A44gBnrqP4OlXFP0pLvcEemdpe7
pg0NoEQC98pwxjGYB04TyUXrCfANUtvbhZFuzQdyA0g0pYdhSg/FAmwJwsJ0stpkWWzPkPNf/GXE
7ZuB329fKYpqgjjZmxA2/t849T82AsmaOLPEPnK/wiSlnvX0hMBbOUW2SGaxkox24yv3loHCiVHr
0kfgEzBcu8+ckSQA7GV7dlq81zGSB3vXhoGYcZVeSe1ytmJwAorHOnuK6KgnF/DOa3O5/w2TVnfF
K5rgWSDgNC6HuvnBX127+P+xoUgbcN3/0A83aTpN3tqAsiAbs8NXKn/LhEm1t2Op/M6KLcT8f3kR
jbQu3711mXnUu8MoQoPCuE+1hlYIC3juat9WKziLP7aqMwyywbij2KSLZ4KR5+a38QoGT392yB2S
i7x7TnwnyzzvEXxQc/H6A/3EyLx6kQ4yVnoG3/TOeucY0Josk2L8ZkychesK0huGtWNLNs5qv2aL
bf0nPPy+Ve1D/Ecl/iAsjNqqblouHnCznPw+VueLCfU9F50apB4KZ8TiOiJTkXanxEH/vif73EqR
rbw8EKyZz/WaiGiwMLNXURixazJbi9bSi3tpC6shu/yt12DvEyggi0Yt885fl9P8R41bavprp7Od
KTTIBoDHAviQu4yHtZjqeBHzRIRkxPqIq4/4L+mmg6w5NZPm3Lqnsto6PxnQD0SRkA/9wwc4fm4W
UfHnQSPpSPnQNFfApD77NlyX5nzUaW6a50EiJjJQHIqNUbQw5jqnQb4PZXdBSvmVqgo7pR0G0bEo
q34oqlvnqaxn1iO9+4ziNicbkEVYhUrdZMdDhW1udGzzRL2Xp6DwTyfMOzWO28K6z06uhdZEBvKU
/zk/rJgdxCaLBoAAMtN20fQC4tgUcfMblIF0hSEUnOwuX+L+p+ZcUPlyc4HntbuTKOE/sVbIcexO
YweXGmw5AjOIzcI4+JGjBWoExuLD7BRJ95Oj/eCrbyX3bEOFgvw9r7X3KB7Rwo5bKWTGU51NxAQ7
RR5Ri3GMZ12whZERCA+mbPT/jp3bEv70ScN5Tkij72rLiMS3YS+kJpneYtNiZvHwv9bmG0qekrJq
dozSlU89EYukubZ2Akt91Ss97OXvo+J3/uznPdNXVQBopS2uYGP94OBBou32rcWDzhTucReKGGm/
5zWT+ouRMc6673la2XSZJ6zluK2ct4DljHQzMrTusofWr5LelPVdI4WXQ7RUtdxD20jYQl2IQjPc
CeOgl2dHU01wYcva6HCB64Qex8kf4KIr4P9Qa8uWRV7r8UBj8pjeqH2MtNwEJ9DbsmmKFdSmp1mN
5x2jcp74ZO8xNEl/wOS0YBIQZilAusXOOediWLxuAAXVy6ZL+M5qFFjSCMO+2kpALztIjvs2zIJA
qnFvwfxY+BesiNgf05e7ORMICiQ6O7uCvb2n9UdQFWVk9+Flv9beD0m6bWOdmMPl0KDYPVO8nlP9
r9D6VNoZHleNvMgQuPFoQap3RxFrIP3WwIdcoCFYGgTWkIiST9Z5FEUluMT4pb7T2qk4f5G3bj9E
HyzuXRyW74m6Qx76z7y/1UnqGnRIkGq9dIZlRYny+HhExeiBzDYQxhiTUf0+TPbtH2HwsCXWLuBC
xJaLtYHqpUBkqdg+BJtqeT13uHlAmx+HxoWgvhJlKXItPsMX/F6Dbi189yyf+mcEp3F2X8TLTXiq
QFjopzKYPzOuD2Sfy+OWgrwlV3Zriw0yrGiTM5TfLN26SBrsBz96VCHQhE4GBMWBgeD5tNB/3wUQ
iQal0qetEuM0kO+4D4sxroflbyZi2+fGP4Utilsy/NLv3HCxZjYb8cuuBgaCvI8d8/x0NfV+d45q
tUTxEdBh9iQnjHvkh4/JONhHLrRFWKFZsNkKkmC48HrX3jXH0ggJt5GBUswJMOU9k01GfmIkJfdE
CLRP4WSBq4RgPw7orHeIt5EFF2c3Jt27LWrrLAMhESgTkRBK+Otg3rMMriHqMh6GeJZOKXasVTEw
qUkDSY9jV7OMd78Y9PmofLjttDcBOskAnWv9NUx6H39Di3ubvHPNDDXT2YgHFvBS8d8JjKzrwLiI
sFhMW+0dG+kdtnfLxDaNXlhw4ul/PvwjQhX3OwwE6YTxJc66c397wRDvkHppQSKtddaXvdGNkT+9
QjTj/qrhkwZ4/LUcp/HTyNHwoPZMX6hsCqhTznSekWJyvXJ5SSf8JHhLIY8i4U6Tt9HfQT5qdqfZ
LXarhKuZGse0u7W5WMXJTcy2Z9ZQONM1SaH9/4r8buTIH3CNi/nskhYLkYOJi5F5lUIcdnHG8EPU
XCd4zZ/0YQV54pb8EJY04aAZhL/EN6W86NUH1ovkWKJrc8FkJQQIKqvqCjQbpDORuiKwkXi9acd0
bx3DLiEUgNLivtwPQXUymmA4EHgbXTU1azvmlaEX2KX4BSMjzlkfsh0S3pH3tacH7Fq/KB39emN+
CmKNuzy8h1XDbGexPLH0csEzn9dEeDsLZNwbBLqIL9n25g5690Bj5O5Vtb7qthUxE8Xs6eUYofFg
1NtDU11snny9FNm29cvbb8MJhiSow07FXwtLPTAOh63ECkcYMvUUp68OZfava1uoEYGuBQkXcxsL
lra3cWkrzMV9SOgYnW3pvqNa1xl5fJYwg1JGGs7dyH3FGY5dNICRA8eYb0e8ehfjA2gpYpKP4hlj
8fzYWDhydBgZVJfQeNZKyIhxLnsE8OFiNlvSXcNny/2Li1Po1jl+6BF7uH08wKbGyE3N17Hh8E7R
o9Ulq9WT/bjka06tNUPu9yjiCURxp4DlqFWVBW4qHkNAPYtVT7MsTIrl+flQNk7nL1zIjhpfmERI
hVot+7ACWNz6mbsULy03itMcudvN5aKtqTp2hSh45QvTOv1Tn41mcI5G5+eGTcW30vxdgLHrg+dK
cz9xF5BVLSWuuh/vGkkh6BYN+HpK8RsYaV8wBwf/jT8ghoqYlw9CX1xbNdOg1Ku0tWq14OxJS/Ld
zj4weot+CVahbsNYH4CmmbK3VsjHVidmtn2DdQwi2Fq+qtn1gw48Qasu+6LZjx51jJApwf4zGGs8
m1uhxVGUbS5fTHcdfc86BnNWMsfiO/gY5EDEruv7+rmzQhjCuFPqcYJHDpGKEhrh4xovGiK+UgLe
hvrxU+vuvhG7bKa+dgjfGK88sxEwv7mMFNBMrK2fGaZX5BlkXtWKXEW5MFY3cPWfBcrlQqmisNMz
zpDW6bJRypMuaL5HuKWWt/2BHr/6wH3CHBQhwip26L/J9L+oR3SMxa5L+NoWVt36yfY47aDB9iPq
pkwuEzmfbgamZjVvEG2aZr8qUz6QksBgAQk6tBzexcuHFtXaZsgof1RXmcaQ/MI5zinZ8P0tgFes
xLi5wDla50rdnYZz+0ZrdhyWJnIcw7BAmTFN71ccH1lpt/MwRZlvn9SnIhZaCbiwHLkSym9GzDge
z/uEL3Bo3TNiqR+iVLzF/LeG5velRIjOnSwVXPcYo95IA82yNZlgpGkAitYvm/QJZsgP6QwknUAP
PtT0zhpz4kD6xtKkH3jwtsb3C4sWPAoGuiHym5+AOHe26r42J6GTQojjPa5Ue2qiNNEU0BJuqMbu
DeTVciwUBL7ifWorV8bGo9ISISr3AD8AzHo7BRZNeJFTlVUoYU1KOULhGcE8d78N9l1d7oXp9xtN
NgW/QhJaOA2134Ea2A670Ox1BT4MA6HTsPGfXxEPq6X6ct+xjn7u9exrLecvZK0xMIPo6zV4QmV9
ZmrZWfp/TAI1mBRdhewcKB7BdCJFxo5fIAt/DsywDTLhsKdfsz5jZuAF8iVpRbWPLjkpyv1fNLij
jYsDhxiGAD5d8pTwFYREYlPfcxcaDp3ZEZr0HPznUdNY3D7ZucxDooyKRbtgC/tFtEkm3E3eQ837
nGucDJYPfpjfGn9zq8OsWrB/6QMpel8xj+j0W/ElRUa2kv18AljoVdTPdxRoJrzY1llLgGMKVSQJ
QxI/990U+YhgAC9rO/L80P6KKlHo+WhF9ww9SO0Rot+6YW3Et5+Hks0opxzrBwZX6euQ6DNmrlWe
3ws8L8lFFL++y73KeXQu1UG7nWm2c4qioNLyM2IEiQfJHGqisO3VXRkT6ZZz42J2FkyYsQHdePaI
o+80lRBwzFMBoS8dJ4rQ5p2IvzNiRwGIVpoRWBA/uLSFntQjqsQxT6QHOaCrq5vpFSOnhGYzVLz7
YMl+v/WcrH6xmRkdWpFWSbpfKSLbCS6SVJDJZqo3zUdzoqtpN53rRtOUzBPno5+j8ykdr3uOmd5s
IHzQkW0VQyshnUUvN0hrsSLsHRgLSj12UFStfHjUbrM/sIfESiuMWNGQAEboqevLczNNmYCg+H7/
zPYujLZjlknrCtQRbQvTcl2ngc5LYgZ0IEkubh/rQWYvHLEIWeE+PLCV5OHtIqqF1UmC2+KgGgMW
r4xdYViOfdmNbpK1tCpmSRYJmAmvFXpQfo/ru/Le5n1++/f1c1v0bGHewgQtuyR9DUa+hSkgfwwx
fUDhYbpknXglT1xz4jQX/RtGvz2C6eFpWIVnSLm94Ru0O/amxhYSdie+GVR+4GqcF4ATKMUFHQJy
TotW9AyqdIZdwGsk21/A0glTKITcUgIcE1vj0FF9HDlogR0qiweoXNcyu93uxSDXA54f4IGUgrVU
flMoEcI/wwEvqPNBHsLKSced6+X/frgOi6KbT0RVNTSa4gIWURwq9D5RTTu4NNw80Pr/NfpMfpDS
HZCeD7PH7YFHYxcRQh830P8G/JUV0AxX7yirpXRCq8YCxKw0myrL92a1DKxIXpqBfXOB44H3EwwV
m03o3J8Xfc2yj49nQrUJw4ngeDPghogsOkHKVfYUhfyI9N+gZcvqq8LITIEt9WYNPjMKygqmEoWy
cs3LGmQIYw6IQPkUz8+VIUBMb6kCdNBFsnRUp/k7mfrRQmH++h+JrjRQtOpsSOKZiYl79cYOkc5h
zGIxwk7IpzOntYy2C2xiH6mjXvMraiH/1FBS0+W7G4KDa9y+WpUmKOmjNzjca+vmRMSeTWmcazU1
EwXkdaA6MONFJfMcXBr43h7cygzEGt+pov2jK+uOAA/lNvnMNMG9tD/1vIcy52XQ2m6yGN1n3XZ/
JJOodJQNa5fm0q7ryOhwXbs/nIJEHmtZi7vTo6u0hJlqivBpw5q/7YQinGwbOfdJYwcZCVRVEcU+
WiURD0/B1R/R9UcaDzYZmGaACv9jW7RWizfvFCuAEDa9oMob5X91hao4hz93S4y7pdSNlNg//BAz
1jjgl7AjcP6rOG61YViOBxCRFtr+71dCHS6U1mHTtcVJWE3IhjUPZx+YIx8yM2bcCCMRUpb/8Wrc
4ssQcUMQX7GF9coJo4sDePgIVq0b9xqga9t4P2luBfs2Q5gOJlBrY+tQnO81HSqaa4gNzKWfUnyQ
LOip2ENTQTcL7EsW+jaDVee08EsN/kfI4IK0zrQ6FneZm5tNNOsgIFMEL4QKvcAV5Uxx8kME7BcQ
ro+kSpdblT2lfZ1hDV0TlSvX8w1laqVUV2dgQ+gYEiPmiFjkz7zQDpX5JQBOWwXRWSkGlA4TNb4e
yDTAc4UzXAsnXGncu6bPTllPeXKd916uy9DpMQngWJ/xtXEDbWrbtmzr67jD0kGe6YG5BOvPT96/
yDoGXvowbHZFhuYDAu4xgHGXhpSRHPLVYMN0B/lwe1XE/psbiucUkmgW096l/9sVUcBcnH9oBYs5
8L2hfwDQvslsI6dOSIRGZ/pOeaNGhwT2apMy8gLVM/7Ma4KNfdJKCBTxF6DeJcfyVuvG3BtaPndk
pbJqivhVSJyUVnXeJQi43vsi1VLnjDofNCOW6AnPXM6Qdpfnz5ssdvxe0gTxF03JynB+GyHJoOb3
QCJFiLu4uCkZjEcvhbah81g2TjBa76DhKTZqZ1E2ENt4ujPpyW6BPZFOMwGW6WDz4tdlyFMfX4C8
PxeRlKlbiPWZAg4ZdnIovvPpy3rC82xTKHSS+4jfWbAs0K5vyWj2X4w8Vs2opg2Dn2sSKR0+Ghn9
6wykOeEGrCeFWrOpNeYyzAX9ZmS7zVWNBsZxwPMtk4uU3K5CGefm05+yTG+Vd8sXpzXRtW8hz6NN
Hw0QnJ9j9HdTlmHKjedOIfbtJfGIS34mvi86t4Pqrvm/NvXjAFQDpZ5JrteVr7FGGzA5VBDTUFO5
i+G+smAzDurXyVRWiRFJKeZtZSR97VBdMsegcKb/in/Z2H8yuT6MRsGJ4xu5C+AStxRGijYP0eR4
6ODbW+NXAStxYjoRPEWOQfh3+3h6R7mWOSFTRIqhvo6/L1lDzS/ck8jxXN1AA0pEalzxNUeC0Crr
PtV4CK5Xe3rJnUiZ598UaMJ8oet3/hGGiqYmnKUN4ZhpswBmFqj0CYsaVE8XNNUYIwP6sbsOwkEC
W4b3qcXqjp0lGR/d/YMsc+AjDPF7wjGiWbG2EcqfpU18wR3GeELdNmmO4UTt1tKv/RLzAYnP5e1X
kNLNnSyU5YY/9uJHPlqe4CZ5KogSyFVibJ8RxDaUa8vSJLKy7dtDM25UxYsGy8KJAXuycM2LRU6W
W+Xl9je79OvD27u2Ndat9/QMgHZsQ5IywUe3sCwpxtXE2Jt6fRxhrQW62ag64w2b0MzJoLJpzPxM
WIsqFyk6IR3DqjjhktjYYWWupYgH+aUyNEZHWJa6lguxsk3TvV8hCpVUDNXXU6FAagpYvhl8qLU5
AEVgctjmxpVUnwkf+bSwMUpDY2R/LEISRere+EVwvDV4jZ9CKlolGsa0RNBawKyGDWYHB5VHeat/
zKSh99yAM7+8N+5ErN0HRDqwA7GSKQLZ7Ga0puHZwBMzitRSaWgbOkp1Cq7VEtTel/C6a9Oands+
EgVlp/zqD//JtfsYYX/7ulnpEAeXp/rDrtRkdWtAmUdTzlsSrXnDx2Loi9TvIZoFpi5bwd+PWm4s
ihdH79+DYa4Vy/nMQn5U5dGUUvHBqrORbpjz1oRrlnYD+JTfT5N5JRHbNTnJESW5O9cbKlvavmSV
aWJGuchwrkyfEp81opLlH4Oz1lR5Qk7erm5y+11j4xduc3+xLVt7tiw9Fc04HzD60EGAnWCYCJn+
xKYtGzxA8NVJZ78GSlbiKq00/0ophtgmsrXqSkzt1MMn67RBZwxdnFQ567u+kl/4LyIE/MB7vLTv
d1qfPjTEAehyw8+VKmVfPr/lvTPzsqa1UWbmjHjCzb0ub92ilhw9+u6q89NVUgAhmNZh/7B4X5Y0
Vtj+/tMz/VpILZi1FXYHU75JVgzrob4N4V39jV6yGEKIfZuuT0BGA3c+IFc49wnShwEZkzmly0o1
SIqx8rTOSUJqcU4tSg4ltCiGZCKb0iQt9CxBtP+7QhaRkwg3CQ9mIWpHkVznhchixBvfauDUzgQE
veul5bizWioOs7z/nYAGW/WUzeSDgzyWf9q/41uqVsufbcDSyWNcSbsnaj5y8BMopySqKTju8sTH
aE5gJYtFR+ZliWhmLoY/NHkNwKYbbfPKqzdIxWbFnVaVIwZfe8+e60Ms+pECSKWUtUrkqbR240ah
7MdHdA6x6/SfIGrakWahPAzUccFxI93n3O5/9O6i6oQfHfr3hHTtXUqZgcAzSCNnEKIyxzV5mvcC
Md2rGaVPAdwQB4t8hT+zq14sPUui9o1x+Nsq1FXjMZ4wtujgL/GNXFjpkHb0jLRd/FA9gMjwTQXi
kElHonyF1atVe7vu5T8SKRDRMpN2U42IdcRsxZhKARhkO0deTVhW3QgLJPTaH0yIHfQb2pGU6Dcy
2Akc8Gj6YWPeNSsnjzqcxs1zzxV2KdjXCNRxDZItgV1X+zzG2hgSO9NxfY1yI2RsEc7KHpJkjZhb
A8Y60BAtgDxEzsk99jhT77v3D1mZFAMzrQYSjhZ1EUvdpBXg/mYVuU1Eqry3n6f6X17AtI4rQUV2
+XGsqExYvC48iw6MUxZegHhu/4CR0+oDUATH0DnM4yu8A8JzufVFSfHMy8ql22JtD2QpbW8BGSRY
tgky5DIdiiba5g7YVzCulWyV469PN/w11YXzysZeMeIrRwZ6iWQvX3TNcb2coTx7jV2s9yZZpuW/
m1p9IxoGufY5M1SCzqZYGC06cvEMzPyuM81pHrJS6b7YAFXBnAr3PIQFc1FbyyYa6b6JVjsYSPW2
CduHpl6RP7wJ3XJ/EUI8XqkuqeVNxtbJE2QhkLSE/+68AZYUEIGRrN8ktx51ButuQFWTJNndgeho
Aray6kdyVVRX5QUUM+i41NLewlGa93M7PQxPX5O/pPIfUQSo5VEauYtOHpx3Pr4lLzST/X7ws1Nq
87oPSDCDRIvvwXvag19KoEjbxmFEh4skvJWL7/yay+fAPlX3JIIgDE9RBtlmXShJIK/xV+nCHgUz
YIaAxbsVmKZ8SK2cEXe9Z8BrDC3QIq35jpxVYuts9H1ToKvzuNWjdgi8HFChZFgV3zFX14RYnqov
gBxKgG5z11PQcYkyD0BQ7qkshnr0e8GYkIb/STaZpCZ7Cr44vlBU6+x9teMpQi/QFbRIGac+5CDt
4ZRlyNWvcnu7Xj62/rQ9S8wiSyc63k6WLoBPHP18KFRO6vcymMD9KTAN9ys6kC696XIm1IWCrUfw
PtVxValSKGlGRBZevbv0kaPrUCnnkK92TDVHt32b+p1jKAX5QtT4aL5G1Aff7y8wKE68wb/Mao+E
L/Yr3uq9MJ7fKwNZOBTTxhy76d8GsHN/J9p+J4Mdp91565YEDxjXhvwDxzsV/xA2OkgFeRyA3l71
/4eHsk2SDq8fUGcyPIyj9Fwzo911S/ofR6AoyPEuTZiaRRlIdSfa5Dwpi9INTzYpgpp8qD8PRBpt
b7xfKhrctZ7ichqn1U+vEeIaMrRMbe0Xze8iZ+SkwaQ8ADB6/355ocicse60hYGgRa80jE6ScKLW
yeIFmnca+gS4fNsq50VSjUlC+fPerZQ8TUMJi5snnlTR1r3NBJKIc8wZsKI0DAUC4sv0Q0wxGROc
wVv7yMPIOJ6YdCs7uLp0rsxShrrLocYgrWvei5Vh/XBLQfFq5pH4Ute3cy4M5Z2ehLksD8uVjXbu
Tcg6sU2E9a5i3WfdJskDZDedhLF1kKqgkcY5/04yWWUEk4bF0rtrUkV8pOXOFv2F61lYZpBOL2vs
P+bKEdP8aF1txhlA8YkJTGW8BSHIDVukxf8FRBPffOVsjr1xpgLKmf/rl5NMQk05slinIoj9Z9Be
Psmqf56lRQTytOGa/2vWsk2ebJ3OcuS13+/KsIV2MIkeAc8OLSN4CQpJ8ZF1pSXAfiSBEditIs6R
Gc/pTVvgTckGnvzTE/z9vUE97H7DdbHimUbI3siX9HV+dpNDUBhcnDVM3ISbGkZcQv3jfdVLZhof
+EPlVofvzNqO47F6lTkHKNOvlhF9q6H5h9hX3o3iawWZc/ZMBva9pQECI7vmoP6xd5TL1FGZMWjd
LLh1N8fOyZe1OWtg93mqEEZjD3/HoVogNaNu0GNMsQ+kQXYTpcnK6RdPJI1J02iKeVv37nf1dfrj
zbvXXi3zgyGCl+OFuf3MK0WIRqHDfOmVNA6HaJBMGyC999R07nawfSuXQ9KnaJrC15KmTutikKlF
lyjaOtHeNPZ9600lmxATAsgu7W79IKbOpbM4PGrcdrqrEA6PZC4Rc+bQ9AY1yhPPLYsLanqgDdpV
u+5hLkCs4iSulddhG7SzgDdTkrRRyYZWk0ueqzkCkf7pt/x5vQUU7H7xtA/lmcDloxaTDezjMXCF
mnLlf6wNfG4/S8/aHyArLGVJS+WvegO8JQzaL4229kQB2CtaiLWGx3j5cCxxJUvDH+F/iAfDrMOK
Ksa2NpnMEuLqE+ZhOEYbwIaIlwVg5Jqz6vWkoZIfbCYAk4rK1ZUWKQG+95Tumrj9cg75O1eWis62
Rx5qAtK8LyI26aZoCC0rWHO71v+YTkTN5tt1ixBjlCvrSIO7aBY+B0LhzjVDLLgqFF7Kn+0jurb6
IuJnF2durR2NAPWKnGtDdqC9Hz41CQvAl4jgobMHF0HpEW6ErhTAfj1mlTg9oWFCsa6yQ/RSYWB/
tEqnfZxRSwYkqjgaOskg6fkx+HMwRkYPb3j1SzYgdBlHEUg1IIHn8f5Vr5cVXL9Jcx3r65sfJofH
BW4TcNLPilIMLNGMl9cg5sFjuiAsRN05oV7KzOmzk5PCt96YD4T/Qaj3Cn1wcs+0u0eFgjYhCtr7
qluYPomrJZSrx5uKsUheUt1Kmsp1o4l47OIEksQP9VAPvBE2Czt9G6uCmYIzPXGKBlOfUnKX/djj
5GrpZradOCI17iR3pYQAsSSuHDkBBA9XTb0uy+ykKLP2zCrCQeJ8SYunnV2xI6KzB64mOHVssynH
F5nCTSyWM1G0qM/C8xtWRvA8Jjt8pqEPgrqOHfz+K3gXwDvJ8rpvFOyYWKXXCUKzQ/Xoh0HcXNil
ZJYin49fLDXS2yomlkZ87rc5W+gI2+Q/5o+sadopIAD8PNxMTohJ+oZVL9GOvzMExmXzdPEkIkHS
XKOAa4Qx0SrpB20cdsP8m/VPWLvZpl7Ewv3dINFUSwgBod00WDD2QwRDSTzkEozW2CinoT/5ZwxL
UFEpqPDmTT0QQtlkZs6hz1deoBLQvoz4IIGfOM0kNDMOt3xtNG3IMJDhwWt8gPNkC4wwRVn8GDyo
hp6D4rft1xaaJrV7qvmv+SVH5Luc/JHwfKLystKZyq3KbiH22P7fixKMURye8rsdbj8UquS0WeqP
pbyUseUGl+cQgkvd5O+0NjjABqRc9AV54W1H3RybzuetH51GhF4mB/dyO9lfHsswASiaFbwuILje
K3yfBd9QOcW1qEjaY7oOhiCORCwjFXC0pXn48oYKJy5q+jmbUv32ssSijpLLXJ8NkjWmYTpD/Icl
EYNziHLpalnlKKVSdb0OTJR7T9tyoXCji5RM7TEwCJRDz5KinPZDHEcOkNS7xEZK2sKuCiwxRSKv
EBa1ELKbFUtbEz4M6ixQpuM2d99VGu86/JtsMYkuJuWldeMQFCMcAedWwptv3GbziNNX2O2x7TCW
+PYG/5a8BqOzJLUp9ATAScuoWNpiQe/+3VhF4jhXibUsmGftBOTkJLslXwzwgGr+dr8sfnV3DmxS
5MF9Qjp+h5jo3k9vL3gTjODQ+C4+FVrex8aRWLTTDvSknuRtVehbsPyjFRqGQreetnlwpX8RcxqZ
JtJRlPZBKmja0vI7iJ+HXO3Hi8u/srK9y6ZrY0g8kdSm/WfxOJAoSVHZtsrdkvmTrss03eaXUhwe
dXOm2iuaQRdMj0J2dDd2wwFl9l+9RlyGgKhHXWaPAxr8ZkMk+KBfav+87csogN9nT2wuN+e8jU5P
LqVAeQFIsaSSYTkEYpIdRIRSx79kScrPvmZslLosU7o0yqnFtDabQvdBawADDtN6AJGUPwoUC0IP
r2tHNe1GSCyagsagbmfNEiqfygggCLY9k5jRugQ5bFaiDtHgNN+fdSox7HKrhkVAI7WO5jI9Yums
tXDvv1FtI5wV2g6IDQHE69xfe0XRQkuQRzCpJXLQg0CFdFSs8gL3qZfLdm0oaq2QtSpdlnQxMlYs
npvYdxaLtiUqgAZq7DbA9xxi82AEZ0PrINaB1mJETaLoh9aqvHZOgK+BC60dZqPeGb1SduzVO5fg
1J07HCON2VE4/n/xitWayjWkl4PbqSYY0vI7xy2wIUy9JnBOxA2PR5rFIPH/OZT+0eYm/kJYitWk
YgPDdc/jH2T/EMESOlzGnGC1iaFANO98xZO3QHsiy/2f557FMLjM0NZ0z9Muat48s9ilbWnNLtss
XK2AgDL3Z6wkkM42LqtlQg357B5yzTm6dK4sT4ReKSaqaPKIhz62jk+GCYxVhsuwgd/UvIT835kC
UpdjR/cG0C/tgvdBzdAAHcKWXCLr2oLVV+MhQ9yb49GIysLEob51HKGLttJIG5ePbXYev1TP+xz8
uYbEzU06ubi5W/pfi/WAjqw8ucyZQkn2sZKDh3L/sP2FPXtZVU1178sVt05zs8y5DRzBwIPiCoHY
dyiQ20JqaOXsFyZKwLvAB9vGhYeOqcS1M0bmGDAYEQ4yBPqMxCxqYrM2bFyGtDIR0q1RygX1h3nM
JWhMCQdh3/lbFwp8y8iJ1DmbrbU0mAV7+EswC6TYJOCXACAZFbZPV0PnYKUQuDEss3F+hcVFU7rk
+NCKpbj4tVFJHeG88AdJtXXGJ3M8uXG0d8AXChZXyLvy50gpF5OIbilIJcz9GNk1T/NCKyWUmz1s
IMZ/ngjc5yJcVSozuRRsPB+iCWG3h4KzlK85FQ5PfRs80RWdx2HYtFsPy7e29g3qbDMtKCef7tXs
1naZro/Gd3wrCtYuX6wI2iKixI95L2pu8vGa/BbVX5i+2dNdzA==
`protect end_protected
